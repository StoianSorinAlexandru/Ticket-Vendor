library	IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_UNSIGNED.all;

entity DEC_12B_4I is
	
	port(
	D:in STD_LOGIC_VECTOR(0 to 11);
	NRU, NRZ, NRS, NRM: out STD_LOGIC_VECTOR(0 to 6));
	
end DEC_12B_4I;

architecture comportamentala of DEC_12B_4I is
														 
	begin
	process(D)									 
	variable B1, B2, B3, B4: STD_LOGIC_VECTOR(0 to 6);
	begin	
		
		case D is	  																	     													
		--0
		when "000000000000" => B1 := "1111110"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--1
		when "000000000001" => B1 := "0110000"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--2
		when "000000000010" => B1 := "1101101"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--3
		when "000000000011" => B1 := "1111001"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--4
		when "000000000100" => B1 := "0110011"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--5
		when "000000000101" => B1 := "1011011"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--6
		when "000000000110" => B1 := "1011111"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--7
		when "000000000111" => B1 := "1110000"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--8
		when "000000001000" => B1 := "1111111"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--9
		when "000000001001" => B1 := "1111011"; B2 := "1111110"; B3 := "1111110"; B4 := "1111110"; 
		--10
		when "000000001010" => B1 := "1111110"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--11
		when "000000001011" => B1 := "0110000"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--12
		when "000000001100" => B1 := "1101101"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--13
		when "000000001101" => B1 := "1111001"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--14
		when "000000001110" => B1 := "0110011"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--15
		when "000000001111" => B1 := "1011011"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--16
		when "000000010000" => B1 := "1011111"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--17
		when "000000010001" => B1 := "1110000"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--18
		when "000000010010" => B1 := "1111111"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--19
		when "000000010011" => B1 := "1111011"; B2 := "0110000"; B3 := "1111110"; B4 := "1111110"; 
		--20
		when "000000010100" => B1 := "1111110"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--21
		when "000000010101" => B1 := "0110000"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--22
		when "000000010110" => B1 := "1101101"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--23
		when "000000010111" => B1 := "1111001"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--24
		when "000000011000" => B1 := "0110011"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--25
		when "000000011001" => B1 := "1011011"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--26
		when "000000011010" => B1 := "1011111"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--27
		when "000000011011" => B1 := "1110000"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--28
		when "000000011100" => B1 := "1111111"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--29
		when "000000011101" => B1 := "1111011"; B2 := "1101101"; B3 := "1111110"; B4 := "1111110"; 
		--30
		when "000000011110" => B1 := "1111110"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--31
		when "000000011111" => B1 := "0110000"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--32
		when "000000100000" => B1 := "1101101"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--33
		when "000000100001" => B1 := "1111001"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--34
		when "000000100010" => B1 := "0110011"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--35
		when "000000100011" => B1 := "1011011"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--36
		when "000000100100" => B1 := "1011111"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--37
		when "000000100101" => B1 := "1110000"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--38
		when "000000100110" => B1 := "1111111"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--39
		when "000000100111" => B1 := "1111011"; B2 := "1111001"; B3 := "1111110"; B4 := "1111110"; 
		--40
		when "000000101000" => B1 := "1111110"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--41
		when "000000101001" => B1 := "0110000"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--42
		when "000000101010" => B1 := "1101101"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--43
		when "000000101011" => B1 := "1111001"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--44
		when "000000101100" => B1 := "0110011"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--45
		when "000000101101" => B1 := "1011011"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--46
		when "000000101110" => B1 := "1011111"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--47
		when "000000101111" => B1 := "1110000"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--48
		when "000000110000" => B1 := "1111111"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--49
		when "000000110001" => B1 := "1111011"; B2 := "0110011"; B3 := "1111110"; B4 := "1111110"; 
		--50
		when "000000110010" => B1 := "1111110"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--51
		when "000000110011" => B1 := "0110000"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--52
		when "000000110100" => B1 := "1101101"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--53
		when "000000110101" => B1 := "1111001"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--54
		when "000000110110" => B1 := "0110011"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--55
		when "000000110111" => B1 := "1011011"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--56
		when "000000111000" => B1 := "1011111"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--57
		when "000000111001" => B1 := "1110000"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--58
		when "000000111010" => B1 := "1111111"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--59
		when "000000111011" => B1 := "1111011"; B2 := "1011011"; B3 := "1111110"; B4 := "1111110"; 
		--60
		when "000000111100" => B1 := "1111110"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--61
		when "000000111101" => B1 := "0110000"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--62
		when "000000111110" => B1 := "1101101"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--63
		when "000000111111" => B1 := "1111001"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--64
		when "000001000000" => B1 := "0110011"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--65
		when "000001000001" => B1 := "1011011"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--66
		when "000001000010" => B1 := "1011111"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--67
		when "000001000011" => B1 := "1110000"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--68
		when "000001000100" => B1 := "1111111"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--69
		when "000001000101" => B1 := "1111011"; B2 := "1011111"; B3 := "1111110"; B4 := "1111110"; 
		--70
		when "000001000110" => B1 := "1111110"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--71
		when "000001000111" => B1 := "0110000"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--72
		when "000001001000" => B1 := "1101101"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--73
		when "000001001001" => B1 := "1111001"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--74
		when "000001001010" => B1 := "0110011"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--75
		when "000001001011" => B1 := "1011011"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--76
		when "000001001100" => B1 := "1011111"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--77
		when "000001001101" => B1 := "1110000"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--78
		when "000001001110" => B1 := "1111111"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--79
		when "000001001111" => B1 := "1111011"; B2 := "1110000"; B3 := "1111110"; B4 := "1111110"; 
		--80
		when "000001010000" => B1 := "1111110"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--81
		when "000001010001" => B1 := "0110000"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--82
		when "000001010010" => B1 := "1101101"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--83
		when "000001010011" => B1 := "1111001"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--84
		when "000001010100" => B1 := "0110011"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--85
		when "000001010101" => B1 := "1011011"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--86
		when "000001010110" => B1 := "1011111"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--87
		when "000001010111" => B1 := "1110000"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--88
		when "000001011000" => B1 := "1111111"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--89
		when "000001011001" => B1 := "1111011"; B2 := "1111111"; B3 := "1111110"; B4 := "1111110"; 
		--90
		when "000001011010" => B1 := "1111110"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--91
		when "000001011011" => B1 := "0110000"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--92
		when "000001011100" => B1 := "1101101"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--93
		when "000001011101" => B1 := "1111001"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--94
		when "000001011110" => B1 := "0110011"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--95
		when "000001011111" => B1 := "1011011"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--96
		when "000001100000" => B1 := "1011111"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--97
		when "000001100001" => B1 := "1110000"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--98
		when "000001100010" => B1 := "1111111"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--99
		when "000001100011" => B1 := "1111011"; B2 := "1111011"; B3 := "1111110"; B4 := "1111110"; 
		--100
		when "000001100100" => B1 := "1111110"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--101
		when "000001100101" => B1 := "0110000"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--102
		when "000001100110" => B1 := "1101101"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--103
		when "000001100111" => B1 := "1111001"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--104
		when "000001101000" => B1 := "0110011"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--105
		when "000001101001" => B1 := "1011011"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--106
		when "000001101010" => B1 := "1011111"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--107
		when "000001101011" => B1 := "1110000"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--108
		when "000001101100" => B1 := "1111111"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--109
		when "000001101101" => B1 := "1111011"; B2 := "1111110"; B3 := "0110000"; B4 := "1111110"; 
		--110
		when "000001101110" => B1 := "1111110"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--111
		when "000001101111" => B1 := "0110000"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--112
		when "000001110000" => B1 := "1101101"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--113
		when "000001110001" => B1 := "1111001"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--114
		when "000001110010" => B1 := "0110011"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--115
		when "000001110011" => B1 := "1011011"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--116
		when "000001110100" => B1 := "1011111"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--117
		when "000001110101" => B1 := "1110000"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--118
		when "000001110110" => B1 := "1111111"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--119
		when "000001110111" => B1 := "1111011"; B2 := "0110000"; B3 := "0110000"; B4 := "1111110"; 
		--120
		when "000001111000" => B1 := "1111110"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--121
		when "000001111001" => B1 := "0110000"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--122
		when "000001111010" => B1 := "1101101"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--123
		when "000001111011" => B1 := "1111001"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--124
		when "000001111100" => B1 := "0110011"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--125
		when "000001111101" => B1 := "1011011"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--126
		when "000001111110" => B1 := "1011111"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--127
		when "000001111111" => B1 := "1110000"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--128
		when "000010000000" => B1 := "1111111"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--129
		when "000010000001" => B1 := "1111011"; B2 := "1101101"; B3 := "0110000"; B4 := "1111110"; 
		--130
		when "000010000010" => B1 := "1111110"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--131
		when "000010000011" => B1 := "0110000"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--132
		when "000010000100" => B1 := "1101101"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--133
		when "000010000101" => B1 := "1111001"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--134
		when "000010000110" => B1 := "0110011"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--135
		when "000010000111" => B1 := "1011011"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--136
		when "000010001000" => B1 := "1011111"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--137
		when "000010001001" => B1 := "1110000"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--138
		when "000010001010" => B1 := "1111111"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--139
		when "000010001011" => B1 := "1111011"; B2 := "1111001"; B3 := "0110000"; B4 := "1111110"; 
		--140
		when "000010001100" => B1 := "1111110"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--141
		when "000010001101" => B1 := "0110000"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--142
		when "000010001110" => B1 := "1101101"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--143
		when "000010001111" => B1 := "1111001"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--144
		when "000010010000" => B1 := "0110011"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--145
		when "000010010001" => B1 := "1011011"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--146
		when "000010010010" => B1 := "1011111"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--147
		when "000010010011" => B1 := "1110000"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--148
		when "000010010100" => B1 := "1111111"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--149
		when "000010010101" => B1 := "1111011"; B2 := "0110011"; B3 := "0110000"; B4 := "1111110"; 
		--150
		when "000010010110" => B1 := "1111110"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--151
		when "000010010111" => B1 := "0110000"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--152
		when "000010011000" => B1 := "1101101"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--153
		when "000010011001" => B1 := "1111001"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--154
		when "000010011010" => B1 := "0110011"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--155
		when "000010011011" => B1 := "1011011"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--156
		when "000010011100" => B1 := "1011111"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--157
		when "000010011101" => B1 := "1110000"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--158
		when "000010011110" => B1 := "1111111"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--159
		when "000010011111" => B1 := "1111011"; B2 := "1011011"; B3 := "0110000"; B4 := "1111110"; 
		--160
		when "000010100000" => B1 := "1111110"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--161
		when "000010100001" => B1 := "0110000"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--162
		when "000010100010" => B1 := "1101101"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--163
		when "000010100011" => B1 := "1111001"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--164
		when "000010100100" => B1 := "0110011"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--165
		when "000010100101" => B1 := "1011011"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--166
		when "000010100110" => B1 := "1011111"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--167
		when "000010100111" => B1 := "1110000"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--168
		when "000010101000" => B1 := "1111111"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--169
		when "000010101001" => B1 := "1111011"; B2 := "1011111"; B3 := "0110000"; B4 := "1111110"; 
		--170
		when "000010101010" => B1 := "1111110"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--171
		when "000010101011" => B1 := "0110000"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--172
		when "000010101100" => B1 := "1101101"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--173
		when "000010101101" => B1 := "1111001"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--174
		when "000010101110" => B1 := "0110011"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--175
		when "000010101111" => B1 := "1011011"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--176
		when "000010110000" => B1 := "1011111"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--177
		when "000010110001" => B1 := "1110000"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--178
		when "000010110010" => B1 := "1111111"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--179
		when "000010110011" => B1 := "1111011"; B2 := "1110000"; B3 := "0110000"; B4 := "1111110"; 
		--180
		when "000010110100" => B1 := "1111110"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--181
		when "000010110101" => B1 := "0110000"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--182
		when "000010110110" => B1 := "1101101"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--183
		when "000010110111" => B1 := "1111001"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--184
		when "000010111000" => B1 := "0110011"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--185
		when "000010111001" => B1 := "1011011"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--186
		when "000010111010" => B1 := "1011111"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--187
		when "000010111011" => B1 := "1110000"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--188
		when "000010111100" => B1 := "1111111"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--189
		when "000010111101" => B1 := "1111011"; B2 := "1111111"; B3 := "0110000"; B4 := "1111110"; 
		--190
		when "000010111110" => B1 := "1111110"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--191
		when "000010111111" => B1 := "0110000"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--192
		when "000011000000" => B1 := "1101101"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--193
		when "000011000001" => B1 := "1111001"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--194
		when "000011000010" => B1 := "0110011"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--195
		when "000011000011" => B1 := "1011011"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--196
		when "000011000100" => B1 := "1011111"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--197
		when "000011000101" => B1 := "1110000"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--198
		when "000011000110" => B1 := "1111111"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--199
		when "000011000111" => B1 := "1111011"; B2 := "1111011"; B3 := "0110000"; B4 := "1111110"; 
		--200
		when "000011001000" => B1 := "1111110"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--201
		when "000011001001" => B1 := "0110000"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--202
		when "000011001010" => B1 := "1101101"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--203
		when "000011001011" => B1 := "1111001"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--204
		when "000011001100" => B1 := "0110011"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--205
		when "000011001101" => B1 := "1011011"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--206
		when "000011001110" => B1 := "1011111"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--207
		when "000011001111" => B1 := "1110000"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--208
		when "000011010000" => B1 := "1111111"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--209
		when "000011010001" => B1 := "1111011"; B2 := "1111110"; B3 := "1101101"; B4 := "1111110"; 
		--210
		when "000011010010" => B1 := "1111110"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--211
		when "000011010011" => B1 := "0110000"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--212
		when "000011010100" => B1 := "1101101"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--213
		when "000011010101" => B1 := "1111001"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--214
		when "000011010110" => B1 := "0110011"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--215
		when "000011010111" => B1 := "1011011"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--216
		when "000011011000" => B1 := "1011111"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--217
		when "000011011001" => B1 := "1110000"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--218
		when "000011011010" => B1 := "1111111"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--219
		when "000011011011" => B1 := "1111011"; B2 := "0110000"; B3 := "1101101"; B4 := "1111110"; 
		--220
		when "000011011100" => B1 := "1111110"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--221
		when "000011011101" => B1 := "0110000"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--222
		when "000011011110" => B1 := "1101101"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--223
		when "000011011111" => B1 := "1111001"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--224
		when "000011100000" => B1 := "0110011"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--225
		when "000011100001" => B1 := "1011011"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--226
		when "000011100010" => B1 := "1011111"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--227
		when "000011100011" => B1 := "1110000"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--228
		when "000011100100" => B1 := "1111111"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--229
		when "000011100101" => B1 := "1111011"; B2 := "1101101"; B3 := "1101101"; B4 := "1111110"; 
		--230
		when "000011100110" => B1 := "1111110"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--231
		when "000011100111" => B1 := "0110000"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--232
		when "000011101000" => B1 := "1101101"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--233
		when "000011101001" => B1 := "1111001"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--234
		when "000011101010" => B1 := "0110011"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--235
		when "000011101011" => B1 := "1011011"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--236
		when "000011101100" => B1 := "1011111"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--237
		when "000011101101" => B1 := "1110000"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--238
		when "000011101110" => B1 := "1111111"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--239
		when "000011101111" => B1 := "1111011"; B2 := "1111001"; B3 := "1101101"; B4 := "1111110"; 
		--240
		when "000011110000" => B1 := "1111110"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--241
		when "000011110001" => B1 := "0110000"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--242
		when "000011110010" => B1 := "1101101"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--243
		when "000011110011" => B1 := "1111001"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--244
		when "000011110100" => B1 := "0110011"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--245
		when "000011110101" => B1 := "1011011"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--246
		when "000011110110" => B1 := "1011111"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--247
		when "000011110111" => B1 := "1110000"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--248
		when "000011111000" => B1 := "1111111"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--249
		when "000011111001" => B1 := "1111011"; B2 := "0110011"; B3 := "1101101"; B4 := "1111110"; 
		--250
		when "000011111010" => B1 := "1111110"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--251
		when "000011111011" => B1 := "0110000"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--252
		when "000011111100" => B1 := "1101101"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--253
		when "000011111101" => B1 := "1111001"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--254
		when "000011111110" => B1 := "0110011"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--255
		when "000011111111" => B1 := "1011011"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--256
		when "000100000000" => B1 := "1011111"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--257
		when "000100000001" => B1 := "1110000"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--258
		when "000100000010" => B1 := "1111111"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--259
		when "000100000011" => B1 := "1111011"; B2 := "1011011"; B3 := "1101101"; B4 := "1111110"; 
		--260
		when "000100000100" => B1 := "1111110"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--261
		when "000100000101" => B1 := "0110000"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--262
		when "000100000110" => B1 := "1101101"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--263
		when "000100000111" => B1 := "1111001"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--264
		when "000100001000" => B1 := "0110011"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--265
		when "000100001001" => B1 := "1011011"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--266
		when "000100001010" => B1 := "1011111"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--267
		when "000100001011" => B1 := "1110000"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--268
		when "000100001100" => B1 := "1111111"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--269
		when "000100001101" => B1 := "1111011"; B2 := "1011111"; B3 := "1101101"; B4 := "1111110"; 
		--270
		when "000100001110" => B1 := "1111110"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--271
		when "000100001111" => B1 := "0110000"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--272
		when "000100010000" => B1 := "1101101"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--273
		when "000100010001" => B1 := "1111001"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--274
		when "000100010010" => B1 := "0110011"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--275
		when "000100010011" => B1 := "1011011"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--276
		when "000100010100" => B1 := "1011111"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--277
		when "000100010101" => B1 := "1110000"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--278
		when "000100010110" => B1 := "1111111"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--279
		when "000100010111" => B1 := "1111011"; B2 := "1110000"; B3 := "1101101"; B4 := "1111110"; 
		--280
		when "000100011000" => B1 := "1111110"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--281
		when "000100011001" => B1 := "0110000"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--282
		when "000100011010" => B1 := "1101101"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--283
		when "000100011011" => B1 := "1111001"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--284
		when "000100011100" => B1 := "0110011"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--285
		when "000100011101" => B1 := "1011011"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--286
		when "000100011110" => B1 := "1011111"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--287
		when "000100011111" => B1 := "1110000"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--288
		when "000100100000" => B1 := "1111111"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--289
		when "000100100001" => B1 := "1111011"; B2 := "1111111"; B3 := "1101101"; B4 := "1111110"; 
		--290
		when "000100100010" => B1 := "1111110"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--291
		when "000100100011" => B1 := "0110000"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--292
		when "000100100100" => B1 := "1101101"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--293
		when "000100100101" => B1 := "1111001"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--294
		when "000100100110" => B1 := "0110011"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--295
		when "000100100111" => B1 := "1011011"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--296
		when "000100101000" => B1 := "1011111"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--297
		when "000100101001" => B1 := "1110000"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--298
		when "000100101010" => B1 := "1111111"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--299
		when "000100101011" => B1 := "1111011"; B2 := "1111011"; B3 := "1101101"; B4 := "1111110"; 
		--300
		when "000100101100" => B1 := "1111110"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--301
		when "000100101101" => B1 := "0110000"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--302
		when "000100101110" => B1 := "1101101"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--303
		when "000100101111" => B1 := "1111001"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--304
		when "000100110000" => B1 := "0110011"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--305
		when "000100110001" => B1 := "1011011"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--306
		when "000100110010" => B1 := "1011111"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--307
		when "000100110011" => B1 := "1110000"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--308
		when "000100110100" => B1 := "1111111"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--309
		when "000100110101" => B1 := "1111011"; B2 := "1111110"; B3 := "1111001"; B4 := "1111110"; 
		--310
		when "000100110110" => B1 := "1111110"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--311
		when "000100110111" => B1 := "0110000"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--312
		when "000100111000" => B1 := "1101101"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--313
		when "000100111001" => B1 := "1111001"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--314
		when "000100111010" => B1 := "0110011"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--315
		when "000100111011" => B1 := "1011011"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--316
		when "000100111100" => B1 := "1011111"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--317
		when "000100111101" => B1 := "1110000"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--318
		when "000100111110" => B1 := "1111111"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--319
		when "000100111111" => B1 := "1111011"; B2 := "0110000"; B3 := "1111001"; B4 := "1111110"; 
		--320
		when "000101000000" => B1 := "1111110"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--321
		when "000101000001" => B1 := "0110000"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--322
		when "000101000010" => B1 := "1101101"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--323
		when "000101000011" => B1 := "1111001"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--324
		when "000101000100" => B1 := "0110011"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--325
		when "000101000101" => B1 := "1011011"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--326
		when "000101000110" => B1 := "1011111"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--327
		when "000101000111" => B1 := "1110000"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--328
		when "000101001000" => B1 := "1111111"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--329
		when "000101001001" => B1 := "1111011"; B2 := "1101101"; B3 := "1111001"; B4 := "1111110"; 
		--330
		when "000101001010" => B1 := "1111110"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--331
		when "000101001011" => B1 := "0110000"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--332
		when "000101001100" => B1 := "1101101"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--333
		when "000101001101" => B1 := "1111001"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--334
		when "000101001110" => B1 := "0110011"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--335
		when "000101001111" => B1 := "1011011"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--336
		when "000101010000" => B1 := "1011111"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--337
		when "000101010001" => B1 := "1110000"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--338
		when "000101010010" => B1 := "1111111"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--339
		when "000101010011" => B1 := "1111011"; B2 := "1111001"; B3 := "1111001"; B4 := "1111110"; 
		--340
		when "000101010100" => B1 := "1111110"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--341
		when "000101010101" => B1 := "0110000"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--342
		when "000101010110" => B1 := "1101101"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--343
		when "000101010111" => B1 := "1111001"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--344
		when "000101011000" => B1 := "0110011"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--345
		when "000101011001" => B1 := "1011011"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--346
		when "000101011010" => B1 := "1011111"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--347
		when "000101011011" => B1 := "1110000"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--348
		when "000101011100" => B1 := "1111111"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--349
		when "000101011101" => B1 := "1111011"; B2 := "0110011"; B3 := "1111001"; B4 := "1111110"; 
		--350
		when "000101011110" => B1 := "1111110"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--351
		when "000101011111" => B1 := "0110000"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--352
		when "000101100000" => B1 := "1101101"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--353
		when "000101100001" => B1 := "1111001"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--354
		when "000101100010" => B1 := "0110011"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--355
		when "000101100011" => B1 := "1011011"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--356
		when "000101100100" => B1 := "1011111"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--357
		when "000101100101" => B1 := "1110000"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--358
		when "000101100110" => B1 := "1111111"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--359
		when "000101100111" => B1 := "1111011"; B2 := "1011011"; B3 := "1111001"; B4 := "1111110"; 
		--360
		when "000101101000" => B1 := "1111110"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--361
		when "000101101001" => B1 := "0110000"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--362
		when "000101101010" => B1 := "1101101"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--363
		when "000101101011" => B1 := "1111001"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--364
		when "000101101100" => B1 := "0110011"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--365
		when "000101101101" => B1 := "1011011"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--366
		when "000101101110" => B1 := "1011111"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--367
		when "000101101111" => B1 := "1110000"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--368
		when "000101110000" => B1 := "1111111"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--369
		when "000101110001" => B1 := "1111011"; B2 := "1011111"; B3 := "1111001"; B4 := "1111110"; 
		--370
		when "000101110010" => B1 := "1111110"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--371
		when "000101110011" => B1 := "0110000"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--372
		when "000101110100" => B1 := "1101101"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--373
		when "000101110101" => B1 := "1111001"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--374
		when "000101110110" => B1 := "0110011"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--375
		when "000101110111" => B1 := "1011011"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--376
		when "000101111000" => B1 := "1011111"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--377
		when "000101111001" => B1 := "1110000"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--378
		when "000101111010" => B1 := "1111111"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--379
		when "000101111011" => B1 := "1111011"; B2 := "1110000"; B3 := "1111001"; B4 := "1111110"; 
		--380
		when "000101111100" => B1 := "1111110"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--381
		when "000101111101" => B1 := "0110000"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--382
		when "000101111110" => B1 := "1101101"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--383
		when "000101111111" => B1 := "1111001"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--384
		when "000110000000" => B1 := "0110011"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--385
		when "000110000001" => B1 := "1011011"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--386
		when "000110000010" => B1 := "1011111"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--387
		when "000110000011" => B1 := "1110000"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--388
		when "000110000100" => B1 := "1111111"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--389
		when "000110000101" => B1 := "1111011"; B2 := "1111111"; B3 := "1111001"; B4 := "1111110"; 
		--390
		when "000110000110" => B1 := "1111110"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--391
		when "000110000111" => B1 := "0110000"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--392
		when "000110001000" => B1 := "1101101"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--393
		when "000110001001" => B1 := "1111001"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--394
		when "000110001010" => B1 := "0110011"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--395
		when "000110001011" => B1 := "1011011"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--396
		when "000110001100" => B1 := "1011111"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--397
		when "000110001101" => B1 := "1110000"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--398
		when "000110001110" => B1 := "1111111"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--399
		when "000110001111" => B1 := "1111011"; B2 := "1111011"; B3 := "1111001"; B4 := "1111110"; 
		--400
		when "000110010000" => B1 := "1111110"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--401
		when "000110010001" => B1 := "0110000"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--402
		when "000110010010" => B1 := "1101101"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--403
		when "000110010011" => B1 := "1111001"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--404
		when "000110010100" => B1 := "0110011"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--405
		when "000110010101" => B1 := "1011011"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--406
		when "000110010110" => B1 := "1011111"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--407
		when "000110010111" => B1 := "1110000"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--408
		when "000110011000" => B1 := "1111111"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--409
		when "000110011001" => B1 := "1111011"; B2 := "1111110"; B3 := "0110011"; B4 := "1111110"; 
		--410
		when "000110011010" => B1 := "1111110"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--411
		when "000110011011" => B1 := "0110000"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--412
		when "000110011100" => B1 := "1101101"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--413
		when "000110011101" => B1 := "1111001"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--414
		when "000110011110" => B1 := "0110011"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--415
		when "000110011111" => B1 := "1011011"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--416
		when "000110100000" => B1 := "1011111"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--417
		when "000110100001" => B1 := "1110000"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--418
		when "000110100010" => B1 := "1111111"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--419
		when "000110100011" => B1 := "1111011"; B2 := "0110000"; B3 := "0110011"; B4 := "1111110"; 
		--420
		when "000110100100" => B1 := "1111110"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--421
		when "000110100101" => B1 := "0110000"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--422
		when "000110100110" => B1 := "1101101"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--423
		when "000110100111" => B1 := "1111001"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--424
		when "000110101000" => B1 := "0110011"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--425
		when "000110101001" => B1 := "1011011"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--426
		when "000110101010" => B1 := "1011111"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--427
		when "000110101011" => B1 := "1110000"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--428
		when "000110101100" => B1 := "1111111"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--429
		when "000110101101" => B1 := "1111011"; B2 := "1101101"; B3 := "0110011"; B4 := "1111110"; 
		--430
		when "000110101110" => B1 := "1111110"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--431
		when "000110101111" => B1 := "0110000"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--432
		when "000110110000" => B1 := "1101101"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--433
		when "000110110001" => B1 := "1111001"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--434
		when "000110110010" => B1 := "0110011"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--435
		when "000110110011" => B1 := "1011011"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--436
		when "000110110100" => B1 := "1011111"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--437
		when "000110110101" => B1 := "1110000"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--438
		when "000110110110" => B1 := "1111111"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--439
		when "000110110111" => B1 := "1111011"; B2 := "1111001"; B3 := "0110011"; B4 := "1111110"; 
		--440
		when "000110111000" => B1 := "1111110"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--441
		when "000110111001" => B1 := "0110000"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--442
		when "000110111010" => B1 := "1101101"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--443
		when "000110111011" => B1 := "1111001"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--444
		when "000110111100" => B1 := "0110011"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--445
		when "000110111101" => B1 := "1011011"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--446
		when "000110111110" => B1 := "1011111"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--447
		when "000110111111" => B1 := "1110000"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--448
		when "000111000000" => B1 := "1111111"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--449
		when "000111000001" => B1 := "1111011"; B2 := "0110011"; B3 := "0110011"; B4 := "1111110"; 
		--450
		when "000111000010" => B1 := "1111110"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--451
		when "000111000011" => B1 := "0110000"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--452
		when "000111000100" => B1 := "1101101"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--453
		when "000111000101" => B1 := "1111001"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--454
		when "000111000110" => B1 := "0110011"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--455
		when "000111000111" => B1 := "1011011"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--456
		when "000111001000" => B1 := "1011111"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--457
		when "000111001001" => B1 := "1110000"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--458
		when "000111001010" => B1 := "1111111"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--459
		when "000111001011" => B1 := "1111011"; B2 := "1011011"; B3 := "0110011"; B4 := "1111110"; 
		--460
		when "000111001100" => B1 := "1111110"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--461
		when "000111001101" => B1 := "0110000"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--462
		when "000111001110" => B1 := "1101101"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--463
		when "000111001111" => B1 := "1111001"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--464
		when "000111010000" => B1 := "0110011"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--465
		when "000111010001" => B1 := "1011011"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--466
		when "000111010010" => B1 := "1011111"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--467
		when "000111010011" => B1 := "1110000"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--468
		when "000111010100" => B1 := "1111111"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--469
		when "000111010101" => B1 := "1111011"; B2 := "1011111"; B3 := "0110011"; B4 := "1111110"; 
		--470
		when "000111010110" => B1 := "1111110"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--471
		when "000111010111" => B1 := "0110000"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--472
		when "000111011000" => B1 := "1101101"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--473
		when "000111011001" => B1 := "1111001"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--474
		when "000111011010" => B1 := "0110011"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--475
		when "000111011011" => B1 := "1011011"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--476
		when "000111011100" => B1 := "1011111"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--477
		when "000111011101" => B1 := "1110000"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--478
		when "000111011110" => B1 := "1111111"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--479
		when "000111011111" => B1 := "1111011"; B2 := "1110000"; B3 := "0110011"; B4 := "1111110"; 
		--480
		when "000111100000" => B1 := "1111110"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--481
		when "000111100001" => B1 := "0110000"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--482
		when "000111100010" => B1 := "1101101"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--483
		when "000111100011" => B1 := "1111001"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--484
		when "000111100100" => B1 := "0110011"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--485
		when "000111100101" => B1 := "1011011"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--486
		when "000111100110" => B1 := "1011111"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--487
		when "000111100111" => B1 := "1110000"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--488
		when "000111101000" => B1 := "1111111"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--489
		when "000111101001" => B1 := "1111011"; B2 := "1111111"; B3 := "0110011"; B4 := "1111110"; 
		--490
		when "000111101010" => B1 := "1111110"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--491
		when "000111101011" => B1 := "0110000"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--492
		when "000111101100" => B1 := "1101101"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--493
		when "000111101101" => B1 := "1111001"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--494
		when "000111101110" => B1 := "0110011"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--495
		when "000111101111" => B1 := "1011011"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--496
		when "000111110000" => B1 := "1011111"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--497
		when "000111110001" => B1 := "1110000"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--498
		when "000111110010" => B1 := "1111111"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--499
		when "000111110011" => B1 := "1111011"; B2 := "1111011"; B3 := "0110011"; B4 := "1111110"; 
		--500
		when "000111110100" => B1 := "1111110"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--501
		when "000111110101" => B1 := "0110000"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--502
		when "000111110110" => B1 := "1101101"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--503
		when "000111110111" => B1 := "1111001"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--504
		when "000111111000" => B1 := "0110011"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--505
		when "000111111001" => B1 := "1011011"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--506
		when "000111111010" => B1 := "1011111"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--507
		when "000111111011" => B1 := "1110000"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--508
		when "000111111100" => B1 := "1111111"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--509
		when "000111111101" => B1 := "1111011"; B2 := "1111110"; B3 := "1011011"; B4 := "1111110"; 
		--510
		when "000111111110" => B1 := "1111110"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--511
		when "000111111111" => B1 := "0110000"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--512
		when "001000000000" => B1 := "1101101"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--513
		when "001000000001" => B1 := "1111001"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--514
		when "001000000010" => B1 := "0110011"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--515
		when "001000000011" => B1 := "1011011"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--516
		when "001000000100" => B1 := "1011111"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--517
		when "001000000101" => B1 := "1110000"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--518
		when "001000000110" => B1 := "1111111"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--519
		when "001000000111" => B1 := "1111011"; B2 := "0110000"; B3 := "1011011"; B4 := "1111110"; 
		--520
		when "001000001000" => B1 := "1111110"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--521
		when "001000001001" => B1 := "0110000"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--522
		when "001000001010" => B1 := "1101101"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--523
		when "001000001011" => B1 := "1111001"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--524
		when "001000001100" => B1 := "0110011"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--525
		when "001000001101" => B1 := "1011011"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--526
		when "001000001110" => B1 := "1011111"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--527
		when "001000001111" => B1 := "1110000"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--528
		when "001000010000" => B1 := "1111111"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--529
		when "001000010001" => B1 := "1111011"; B2 := "1101101"; B3 := "1011011"; B4 := "1111110"; 
		--530
		when "001000010010" => B1 := "1111110"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--531
		when "001000010011" => B1 := "0110000"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--532
		when "001000010100" => B1 := "1101101"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--533
		when "001000010101" => B1 := "1111001"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--534
		when "001000010110" => B1 := "0110011"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--535
		when "001000010111" => B1 := "1011011"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--536
		when "001000011000" => B1 := "1011111"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--537
		when "001000011001" => B1 := "1110000"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--538
		when "001000011010" => B1 := "1111111"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--539
		when "001000011011" => B1 := "1111011"; B2 := "1111001"; B3 := "1011011"; B4 := "1111110"; 
		--540
		when "001000011100" => B1 := "1111110"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--541
		when "001000011101" => B1 := "0110000"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--542
		when "001000011110" => B1 := "1101101"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--543
		when "001000011111" => B1 := "1111001"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--544
		when "001000100000" => B1 := "0110011"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--545
		when "001000100001" => B1 := "1011011"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--546
		when "001000100010" => B1 := "1011111"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--547
		when "001000100011" => B1 := "1110000"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--548
		when "001000100100" => B1 := "1111111"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--549
		when "001000100101" => B1 := "1111011"; B2 := "0110011"; B3 := "1011011"; B4 := "1111110"; 
		--550
		when "001000100110" => B1 := "1111110"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--551
		when "001000100111" => B1 := "0110000"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--552
		when "001000101000" => B1 := "1101101"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--553
		when "001000101001" => B1 := "1111001"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--554
		when "001000101010" => B1 := "0110011"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--555
		when "001000101011" => B1 := "1011011"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--556
		when "001000101100" => B1 := "1011111"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--557
		when "001000101101" => B1 := "1110000"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--558
		when "001000101110" => B1 := "1111111"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--559
		when "001000101111" => B1 := "1111011"; B2 := "1011011"; B3 := "1011011"; B4 := "1111110"; 
		--560
		when "001000110000" => B1 := "1111110"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--561
		when "001000110001" => B1 := "0110000"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--562
		when "001000110010" => B1 := "1101101"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--563
		when "001000110011" => B1 := "1111001"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--564
		when "001000110100" => B1 := "0110011"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--565
		when "001000110101" => B1 := "1011011"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--566
		when "001000110110" => B1 := "1011111"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--567
		when "001000110111" => B1 := "1110000"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--568
		when "001000111000" => B1 := "1111111"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--569
		when "001000111001" => B1 := "1111011"; B2 := "1011111"; B3 := "1011011"; B4 := "1111110"; 
		--570
		when "001000111010" => B1 := "1111110"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--571
		when "001000111011" => B1 := "0110000"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--572
		when "001000111100" => B1 := "1101101"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--573
		when "001000111101" => B1 := "1111001"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--574
		when "001000111110" => B1 := "0110011"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--575
		when "001000111111" => B1 := "1011011"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--576
		when "001001000000" => B1 := "1011111"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--577
		when "001001000001" => B1 := "1110000"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--578
		when "001001000010" => B1 := "1111111"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--579
		when "001001000011" => B1 := "1111011"; B2 := "1110000"; B3 := "1011011"; B4 := "1111110"; 
		--580
		when "001001000100" => B1 := "1111110"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--581
		when "001001000101" => B1 := "0110000"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--582
		when "001001000110" => B1 := "1101101"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--583
		when "001001000111" => B1 := "1111001"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--584
		when "001001001000" => B1 := "0110011"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--585
		when "001001001001" => B1 := "1011011"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--586
		when "001001001010" => B1 := "1011111"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--587
		when "001001001011" => B1 := "1110000"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--588
		when "001001001100" => B1 := "1111111"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--589
		when "001001001101" => B1 := "1111011"; B2 := "1111111"; B3 := "1011011"; B4 := "1111110"; 
		--590
		when "001001001110" => B1 := "1111110"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--591
		when "001001001111" => B1 := "0110000"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--592
		when "001001010000" => B1 := "1101101"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--593
		when "001001010001" => B1 := "1111001"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--594
		when "001001010010" => B1 := "0110011"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--595
		when "001001010011" => B1 := "1011011"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--596
		when "001001010100" => B1 := "1011111"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--597
		when "001001010101" => B1 := "1110000"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--598
		when "001001010110" => B1 := "1111111"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--599
		when "001001010111" => B1 := "1111011"; B2 := "1111011"; B3 := "1011011"; B4 := "1111110"; 
		--600
		when "001001011000" => B1 := "1111110"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--601
		when "001001011001" => B1 := "0110000"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--602
		when "001001011010" => B1 := "1101101"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--603
		when "001001011011" => B1 := "1111001"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--604
		when "001001011100" => B1 := "0110011"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--605
		when "001001011101" => B1 := "1011011"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--606
		when "001001011110" => B1 := "1011111"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--607
		when "001001011111" => B1 := "1110000"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--608
		when "001001100000" => B1 := "1111111"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--609
		when "001001100001" => B1 := "1111011"; B2 := "1111110"; B3 := "1011111"; B4 := "1111110"; 
		--610
		when "001001100010" => B1 := "1111110"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--611
		when "001001100011" => B1 := "0110000"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--612
		when "001001100100" => B1 := "1101101"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--613
		when "001001100101" => B1 := "1111001"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--614
		when "001001100110" => B1 := "0110011"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--615
		when "001001100111" => B1 := "1011011"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--616
		when "001001101000" => B1 := "1011111"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--617
		when "001001101001" => B1 := "1110000"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--618
		when "001001101010" => B1 := "1111111"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--619
		when "001001101011" => B1 := "1111011"; B2 := "0110000"; B3 := "1011111"; B4 := "1111110"; 
		--620
		when "001001101100" => B1 := "1111110"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--621
		when "001001101101" => B1 := "0110000"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--622
		when "001001101110" => B1 := "1101101"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--623
		when "001001101111" => B1 := "1111001"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--624
		when "001001110000" => B1 := "0110011"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--625
		when "001001110001" => B1 := "1011011"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--626
		when "001001110010" => B1 := "1011111"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--627
		when "001001110011" => B1 := "1110000"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--628
		when "001001110100" => B1 := "1111111"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--629
		when "001001110101" => B1 := "1111011"; B2 := "1101101"; B3 := "1011111"; B4 := "1111110"; 
		--630
		when "001001110110" => B1 := "1111110"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--631
		when "001001110111" => B1 := "0110000"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--632
		when "001001111000" => B1 := "1101101"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--633
		when "001001111001" => B1 := "1111001"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--634
		when "001001111010" => B1 := "0110011"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--635
		when "001001111011" => B1 := "1011011"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--636
		when "001001111100" => B1 := "1011111"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--637
		when "001001111101" => B1 := "1110000"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--638
		when "001001111110" => B1 := "1111111"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--639
		when "001001111111" => B1 := "1111011"; B2 := "1111001"; B3 := "1011111"; B4 := "1111110"; 
		--640
		when "001010000000" => B1 := "1111110"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--641
		when "001010000001" => B1 := "0110000"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--642
		when "001010000010" => B1 := "1101101"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--643
		when "001010000011" => B1 := "1111001"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--644
		when "001010000100" => B1 := "0110011"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--645
		when "001010000101" => B1 := "1011011"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--646
		when "001010000110" => B1 := "1011111"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--647
		when "001010000111" => B1 := "1110000"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--648
		when "001010001000" => B1 := "1111111"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--649
		when "001010001001" => B1 := "1111011"; B2 := "0110011"; B3 := "1011111"; B4 := "1111110"; 
		--650
		when "001010001010" => B1 := "1111110"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--651
		when "001010001011" => B1 := "0110000"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--652
		when "001010001100" => B1 := "1101101"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--653
		when "001010001101" => B1 := "1111001"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--654
		when "001010001110" => B1 := "0110011"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--655
		when "001010001111" => B1 := "1011011"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--656
		when "001010010000" => B1 := "1011111"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--657
		when "001010010001" => B1 := "1110000"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--658
		when "001010010010" => B1 := "1111111"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--659
		when "001010010011" => B1 := "1111011"; B2 := "1011011"; B3 := "1011111"; B4 := "1111110"; 
		--660
		when "001010010100" => B1 := "1111110"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--661
		when "001010010101" => B1 := "0110000"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--662
		when "001010010110" => B1 := "1101101"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--663
		when "001010010111" => B1 := "1111001"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--664
		when "001010011000" => B1 := "0110011"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--665
		when "001010011001" => B1 := "1011011"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--666
		when "001010011010" => B1 := "1011111"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--667
		when "001010011011" => B1 := "1110000"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--668
		when "001010011100" => B1 := "1111111"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--669
		when "001010011101" => B1 := "1111011"; B2 := "1011111"; B3 := "1011111"; B4 := "1111110"; 
		--670
		when "001010011110" => B1 := "1111110"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--671
		when "001010011111" => B1 := "0110000"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--672
		when "001010100000" => B1 := "1101101"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--673
		when "001010100001" => B1 := "1111001"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--674
		when "001010100010" => B1 := "0110011"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--675
		when "001010100011" => B1 := "1011011"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--676
		when "001010100100" => B1 := "1011111"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--677
		when "001010100101" => B1 := "1110000"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--678
		when "001010100110" => B1 := "1111111"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--679
		when "001010100111" => B1 := "1111011"; B2 := "1110000"; B3 := "1011111"; B4 := "1111110"; 
		--680
		when "001010101000" => B1 := "1111110"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--681
		when "001010101001" => B1 := "0110000"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--682
		when "001010101010" => B1 := "1101101"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--683
		when "001010101011" => B1 := "1111001"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--684
		when "001010101100" => B1 := "0110011"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--685
		when "001010101101" => B1 := "1011011"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--686
		when "001010101110" => B1 := "1011111"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--687
		when "001010101111" => B1 := "1110000"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--688
		when "001010110000" => B1 := "1111111"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--689
		when "001010110001" => B1 := "1111011"; B2 := "1111111"; B3 := "1011111"; B4 := "1111110"; 
		--690
		when "001010110010" => B1 := "1111110"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--691
		when "001010110011" => B1 := "0110000"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--692
		when "001010110100" => B1 := "1101101"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--693
		when "001010110101" => B1 := "1111001"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--694
		when "001010110110" => B1 := "0110011"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--695
		when "001010110111" => B1 := "1011011"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--696
		when "001010111000" => B1 := "1011111"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--697
		when "001010111001" => B1 := "1110000"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--698
		when "001010111010" => B1 := "1111111"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--699
		when "001010111011" => B1 := "1111011"; B2 := "1111011"; B3 := "1011111"; B4 := "1111110"; 
		--700
		when "001010111100" => B1 := "1111110"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--701
		when "001010111101" => B1 := "0110000"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--702
		when "001010111110" => B1 := "1101101"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--703
		when "001010111111" => B1 := "1111001"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--704
		when "001011000000" => B1 := "0110011"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--705
		when "001011000001" => B1 := "1011011"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--706
		when "001011000010" => B1 := "1011111"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--707
		when "001011000011" => B1 := "1110000"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--708
		when "001011000100" => B1 := "1111111"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--709
		when "001011000101" => B1 := "1111011"; B2 := "1111110"; B3 := "1110000"; B4 := "1111110"; 
		--710
		when "001011000110" => B1 := "1111110"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--711
		when "001011000111" => B1 := "0110000"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--712
		when "001011001000" => B1 := "1101101"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--713
		when "001011001001" => B1 := "1111001"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--714
		when "001011001010" => B1 := "0110011"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--715
		when "001011001011" => B1 := "1011011"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--716
		when "001011001100" => B1 := "1011111"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--717
		when "001011001101" => B1 := "1110000"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--718
		when "001011001110" => B1 := "1111111"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--719
		when "001011001111" => B1 := "1111011"; B2 := "0110000"; B3 := "1110000"; B4 := "1111110"; 
		--720
		when "001011010000" => B1 := "1111110"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--721
		when "001011010001" => B1 := "0110000"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--722
		when "001011010010" => B1 := "1101101"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--723
		when "001011010011" => B1 := "1111001"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--724
		when "001011010100" => B1 := "0110011"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--725
		when "001011010101" => B1 := "1011011"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--726
		when "001011010110" => B1 := "1011111"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--727
		when "001011010111" => B1 := "1110000"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--728
		when "001011011000" => B1 := "1111111"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--729
		when "001011011001" => B1 := "1111011"; B2 := "1101101"; B3 := "1110000"; B4 := "1111110"; 
		--730
		when "001011011010" => B1 := "1111110"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--731
		when "001011011011" => B1 := "0110000"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--732
		when "001011011100" => B1 := "1101101"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--733
		when "001011011101" => B1 := "1111001"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--734
		when "001011011110" => B1 := "0110011"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--735
		when "001011011111" => B1 := "1011011"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--736
		when "001011100000" => B1 := "1011111"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--737
		when "001011100001" => B1 := "1110000"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--738
		when "001011100010" => B1 := "1111111"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--739
		when "001011100011" => B1 := "1111011"; B2 := "1111001"; B3 := "1110000"; B4 := "1111110"; 
		--740
		when "001011100100" => B1 := "1111110"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--741
		when "001011100101" => B1 := "0110000"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--742
		when "001011100110" => B1 := "1101101"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--743
		when "001011100111" => B1 := "1111001"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--744
		when "001011101000" => B1 := "0110011"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--745
		when "001011101001" => B1 := "1011011"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--746
		when "001011101010" => B1 := "1011111"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--747
		when "001011101011" => B1 := "1110000"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--748
		when "001011101100" => B1 := "1111111"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--749
		when "001011101101" => B1 := "1111011"; B2 := "0110011"; B3 := "1110000"; B4 := "1111110"; 
		--750
		when "001011101110" => B1 := "1111110"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--751
		when "001011101111" => B1 := "0110000"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--752
		when "001011110000" => B1 := "1101101"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--753
		when "001011110001" => B1 := "1111001"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--754
		when "001011110010" => B1 := "0110011"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--755
		when "001011110011" => B1 := "1011011"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--756
		when "001011110100" => B1 := "1011111"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--757
		when "001011110101" => B1 := "1110000"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--758
		when "001011110110" => B1 := "1111111"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--759
		when "001011110111" => B1 := "1111011"; B2 := "1011011"; B3 := "1110000"; B4 := "1111110"; 
		--760
		when "001011111000" => B1 := "1111110"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--761
		when "001011111001" => B1 := "0110000"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--762
		when "001011111010" => B1 := "1101101"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--763
		when "001011111011" => B1 := "1111001"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--764
		when "001011111100" => B1 := "0110011"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--765
		when "001011111101" => B1 := "1011011"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--766
		when "001011111110" => B1 := "1011111"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--767
		when "001011111111" => B1 := "1110000"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--768
		when "001100000000" => B1 := "1111111"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--769
		when "001100000001" => B1 := "1111011"; B2 := "1011111"; B3 := "1110000"; B4 := "1111110"; 
		--770
		when "001100000010" => B1 := "1111110"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--771
		when "001100000011" => B1 := "0110000"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--772
		when "001100000100" => B1 := "1101101"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--773
		when "001100000101" => B1 := "1111001"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--774
		when "001100000110" => B1 := "0110011"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--775
		when "001100000111" => B1 := "1011011"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--776
		when "001100001000" => B1 := "1011111"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--777
		when "001100001001" => B1 := "1110000"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--778
		when "001100001010" => B1 := "1111111"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--779
		when "001100001011" => B1 := "1111011"; B2 := "1110000"; B3 := "1110000"; B4 := "1111110"; 
		--780
		when "001100001100" => B1 := "1111110"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--781
		when "001100001101" => B1 := "0110000"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--782
		when "001100001110" => B1 := "1101101"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--783
		when "001100001111" => B1 := "1111001"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--784
		when "001100010000" => B1 := "0110011"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--785
		when "001100010001" => B1 := "1011011"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--786
		when "001100010010" => B1 := "1011111"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--787
		when "001100010011" => B1 := "1110000"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--788
		when "001100010100" => B1 := "1111111"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--789
		when "001100010101" => B1 := "1111011"; B2 := "1111111"; B3 := "1110000"; B4 := "1111110"; 
		--790
		when "001100010110" => B1 := "1111110"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--791
		when "001100010111" => B1 := "0110000"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--792
		when "001100011000" => B1 := "1101101"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--793
		when "001100011001" => B1 := "1111001"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--794
		when "001100011010" => B1 := "0110011"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--795
		when "001100011011" => B1 := "1011011"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--796
		when "001100011100" => B1 := "1011111"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--797
		when "001100011101" => B1 := "1110000"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--798
		when "001100011110" => B1 := "1111111"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--799
		when "001100011111" => B1 := "1111011"; B2 := "1111011"; B3 := "1110000"; B4 := "1111110"; 
		--800
		when "001100100000" => B1 := "1111110"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--801
		when "001100100001" => B1 := "0110000"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--802
		when "001100100010" => B1 := "1101101"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--803
		when "001100100011" => B1 := "1111001"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--804
		when "001100100100" => B1 := "0110011"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--805
		when "001100100101" => B1 := "1011011"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--806
		when "001100100110" => B1 := "1011111"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--807
		when "001100100111" => B1 := "1110000"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--808
		when "001100101000" => B1 := "1111111"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--809
		when "001100101001" => B1 := "1111011"; B2 := "1111110"; B3 := "1111111"; B4 := "1111110"; 
		--810
		when "001100101010" => B1 := "1111110"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--811
		when "001100101011" => B1 := "0110000"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--812
		when "001100101100" => B1 := "1101101"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--813
		when "001100101101" => B1 := "1111001"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--814
		when "001100101110" => B1 := "0110011"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--815
		when "001100101111" => B1 := "1011011"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--816
		when "001100110000" => B1 := "1011111"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--817
		when "001100110001" => B1 := "1110000"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--818
		when "001100110010" => B1 := "1111111"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--819
		when "001100110011" => B1 := "1111011"; B2 := "0110000"; B3 := "1111111"; B4 := "1111110"; 
		--820
		when "001100110100" => B1 := "1111110"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--821
		when "001100110101" => B1 := "0110000"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--822
		when "001100110110" => B1 := "1101101"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--823
		when "001100110111" => B1 := "1111001"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--824
		when "001100111000" => B1 := "0110011"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--825
		when "001100111001" => B1 := "1011011"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--826
		when "001100111010" => B1 := "1011111"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--827
		when "001100111011" => B1 := "1110000"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--828
		when "001100111100" => B1 := "1111111"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--829
		when "001100111101" => B1 := "1111011"; B2 := "1101101"; B3 := "1111111"; B4 := "1111110"; 
		--830
		when "001100111110" => B1 := "1111110"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--831
		when "001100111111" => B1 := "0110000"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--832
		when "001101000000" => B1 := "1101101"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--833
		when "001101000001" => B1 := "1111001"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--834
		when "001101000010" => B1 := "0110011"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--835
		when "001101000011" => B1 := "1011011"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--836
		when "001101000100" => B1 := "1011111"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--837
		when "001101000101" => B1 := "1110000"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--838
		when "001101000110" => B1 := "1111111"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--839
		when "001101000111" => B1 := "1111011"; B2 := "1111001"; B3 := "1111111"; B4 := "1111110"; 
		--840
		when "001101001000" => B1 := "1111110"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--841
		when "001101001001" => B1 := "0110000"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--842
		when "001101001010" => B1 := "1101101"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--843
		when "001101001011" => B1 := "1111001"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--844
		when "001101001100" => B1 := "0110011"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--845
		when "001101001101" => B1 := "1011011"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--846
		when "001101001110" => B1 := "1011111"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--847
		when "001101001111" => B1 := "1110000"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--848
		when "001101010000" => B1 := "1111111"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--849
		when "001101010001" => B1 := "1111011"; B2 := "0110011"; B3 := "1111111"; B4 := "1111110"; 
		--850
		when "001101010010" => B1 := "1111110"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--851
		when "001101010011" => B1 := "0110000"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--852
		when "001101010100" => B1 := "1101101"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--853
		when "001101010101" => B1 := "1111001"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--854
		when "001101010110" => B1 := "0110011"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--855
		when "001101010111" => B1 := "1011011"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--856
		when "001101011000" => B1 := "1011111"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--857
		when "001101011001" => B1 := "1110000"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--858
		when "001101011010" => B1 := "1111111"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--859
		when "001101011011" => B1 := "1111011"; B2 := "1011011"; B3 := "1111111"; B4 := "1111110"; 
		--860
		when "001101011100" => B1 := "1111110"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--861
		when "001101011101" => B1 := "0110000"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--862
		when "001101011110" => B1 := "1101101"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--863
		when "001101011111" => B1 := "1111001"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--864
		when "001101100000" => B1 := "0110011"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--865
		when "001101100001" => B1 := "1011011"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--866
		when "001101100010" => B1 := "1011111"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--867
		when "001101100011" => B1 := "1110000"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--868
		when "001101100100" => B1 := "1111111"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--869
		when "001101100101" => B1 := "1111011"; B2 := "1011111"; B3 := "1111111"; B4 := "1111110"; 
		--870
		when "001101100110" => B1 := "1111110"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--871
		when "001101100111" => B1 := "0110000"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--872
		when "001101101000" => B1 := "1101101"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--873
		when "001101101001" => B1 := "1111001"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--874
		when "001101101010" => B1 := "0110011"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--875
		when "001101101011" => B1 := "1011011"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--876
		when "001101101100" => B1 := "1011111"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--877
		when "001101101101" => B1 := "1110000"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--878
		when "001101101110" => B1 := "1111111"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--879
		when "001101101111" => B1 := "1111011"; B2 := "1110000"; B3 := "1111111"; B4 := "1111110"; 
		--880
		when "001101110000" => B1 := "1111110"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--881
		when "001101110001" => B1 := "0110000"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--882
		when "001101110010" => B1 := "1101101"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--883
		when "001101110011" => B1 := "1111001"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--884
		when "001101110100" => B1 := "0110011"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--885
		when "001101110101" => B1 := "1011011"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--886
		when "001101110110" => B1 := "1011111"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--887
		when "001101110111" => B1 := "1110000"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--888
		when "001101111000" => B1 := "1111111"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--889
		when "001101111001" => B1 := "1111011"; B2 := "1111111"; B3 := "1111111"; B4 := "1111110"; 
		--890
		when "001101111010" => B1 := "1111110"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--891
		when "001101111011" => B1 := "0110000"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--892
		when "001101111100" => B1 := "1101101"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--893
		when "001101111101" => B1 := "1111001"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--894
		when "001101111110" => B1 := "0110011"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--895
		when "001101111111" => B1 := "1011011"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--896
		when "001110000000" => B1 := "1011111"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--897
		when "001110000001" => B1 := "1110000"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--898
		when "001110000010" => B1 := "1111111"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--899
		when "001110000011" => B1 := "1111011"; B2 := "1111011"; B3 := "1111111"; B4 := "1111110"; 
		--900
		when "001110000100" => B1 := "1111110"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--901
		when "001110000101" => B1 := "0110000"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--902
		when "001110000110" => B1 := "1101101"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--903
		when "001110000111" => B1 := "1111001"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--904
		when "001110001000" => B1 := "0110011"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--905
		when "001110001001" => B1 := "1011011"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--906
		when "001110001010" => B1 := "1011111"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--907
		when "001110001011" => B1 := "1110000"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--908
		when "001110001100" => B1 := "1111111"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--909
		when "001110001101" => B1 := "1111011"; B2 := "1111110"; B3 := "1111011"; B4 := "1111110"; 
		--910
		when "001110001110" => B1 := "1111110"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--911
		when "001110001111" => B1 := "0110000"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--912
		when "001110010000" => B1 := "1101101"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--913
		when "001110010001" => B1 := "1111001"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--914
		when "001110010010" => B1 := "0110011"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--915
		when "001110010011" => B1 := "1011011"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--916
		when "001110010100" => B1 := "1011111"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--917
		when "001110010101" => B1 := "1110000"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--918
		when "001110010110" => B1 := "1111111"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--919
		when "001110010111" => B1 := "1111011"; B2 := "0110000"; B3 := "1111011"; B4 := "1111110"; 
		--920
		when "001110011000" => B1 := "1111110"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--921
		when "001110011001" => B1 := "0110000"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--922
		when "001110011010" => B1 := "1101101"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--923
		when "001110011011" => B1 := "1111001"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--924
		when "001110011100" => B1 := "0110011"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--925
		when "001110011101" => B1 := "1011011"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--926
		when "001110011110" => B1 := "1011111"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--927
		when "001110011111" => B1 := "1110000"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--928
		when "001110100000" => B1 := "1111111"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--929
		when "001110100001" => B1 := "1111011"; B2 := "1101101"; B3 := "1111011"; B4 := "1111110"; 
		--930
		when "001110100010" => B1 := "1111110"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--931
		when "001110100011" => B1 := "0110000"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--932
		when "001110100100" => B1 := "1101101"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--933
		when "001110100101" => B1 := "1111001"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--934
		when "001110100110" => B1 := "0110011"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--935
		when "001110100111" => B1 := "1011011"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--936
		when "001110101000" => B1 := "1011111"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--937
		when "001110101001" => B1 := "1110000"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--938
		when "001110101010" => B1 := "1111111"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--939
		when "001110101011" => B1 := "1111011"; B2 := "1111001"; B3 := "1111011"; B4 := "1111110"; 
		--940
		when "001110101100" => B1 := "1111110"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--941
		when "001110101101" => B1 := "0110000"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--942
		when "001110101110" => B1 := "1101101"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--943
		when "001110101111" => B1 := "1111001"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--944
		when "001110110000" => B1 := "0110011"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--945
		when "001110110001" => B1 := "1011011"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--946
		when "001110110010" => B1 := "1011111"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--947
		when "001110110011" => B1 := "1110000"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--948
		when "001110110100" => B1 := "1111111"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--949
		when "001110110101" => B1 := "1111011"; B2 := "0110011"; B3 := "1111011"; B4 := "1111110"; 
		--950
		when "001110110110" => B1 := "1111110"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--951
		when "001110110111" => B1 := "0110000"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--952
		when "001110111000" => B1 := "1101101"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--953
		when "001110111001" => B1 := "1111001"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--954
		when "001110111010" => B1 := "0110011"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--955
		when "001110111011" => B1 := "1011011"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--956
		when "001110111100" => B1 := "1011111"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--957
		when "001110111101" => B1 := "1110000"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--958
		when "001110111110" => B1 := "1111111"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--959
		when "001110111111" => B1 := "1111011"; B2 := "1011011"; B3 := "1111011"; B4 := "1111110"; 
		--960
		when "001111000000" => B1 := "1111110"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--961
		when "001111000001" => B1 := "0110000"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--962
		when "001111000010" => B1 := "1101101"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--963
		when "001111000011" => B1 := "1111001"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--964
		when "001111000100" => B1 := "0110011"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--965
		when "001111000101" => B1 := "1011011"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--966
		when "001111000110" => B1 := "1011111"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--967
		when "001111000111" => B1 := "1110000"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--968
		when "001111001000" => B1 := "1111111"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--969
		when "001111001001" => B1 := "1111011"; B2 := "1011111"; B3 := "1111011"; B4 := "1111110"; 
		--970
		when "001111001010" => B1 := "1111110"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--971
		when "001111001011" => B1 := "0110000"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--972
		when "001111001100" => B1 := "1101101"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--973
		when "001111001101" => B1 := "1111001"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--974
		when "001111001110" => B1 := "0110011"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--975
		when "001111001111" => B1 := "1011011"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--976
		when "001111010000" => B1 := "1011111"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--977
		when "001111010001" => B1 := "1110000"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--978
		when "001111010010" => B1 := "1111111"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--979
		when "001111010011" => B1 := "1111011"; B2 := "1110000"; B3 := "1111011"; B4 := "1111110"; 
		--980
		when "001111010100" => B1 := "1111110"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--981
		when "001111010101" => B1 := "0110000"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--982
		when "001111010110" => B1 := "1101101"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--983
		when "001111010111" => B1 := "1111001"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--984
		when "001111011000" => B1 := "0110011"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--985
		when "001111011001" => B1 := "1011011"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--986
		when "001111011010" => B1 := "1011111"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--987
		when "001111011011" => B1 := "1110000"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--988
		when "001111011100" => B1 := "1111111"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--989
		when "001111011101" => B1 := "1111011"; B2 := "1111111"; B3 := "1111011"; B4 := "1111110"; 
		--990
		when "001111011110" => B1 := "1111110"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--991
		when "001111011111" => B1 := "0110000"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--992
		when "001111100000" => B1 := "1101101"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--993
		when "001111100001" => B1 := "1111001"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--994
		when "001111100010" => B1 := "0110011"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--995
		when "001111100011" => B1 := "1011011"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--996
		when "001111100100" => B1 := "1011111"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--997
		when "001111100101" => B1 := "1110000"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--998
		when "001111100110" => B1 := "1111111"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--999
		when "001111100111" => B1 := "1111011"; B2 := "1111011"; B3 := "1111011"; B4 := "1111110"; 
		--1000
		when "001111101000" => B1 := "1111110"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1001
		when "001111101001" => B1 := "0110000"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1002
		when "001111101010" => B1 := "1101101"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1003
		when "001111101011" => B1 := "1111001"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1004
		when "001111101100" => B1 := "0110011"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1005
		when "001111101101" => B1 := "1011011"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1006
		when "001111101110" => B1 := "1011111"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1007
		when "001111101111" => B1 := "1110000"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1008
		when "001111110000" => B1 := "1111111"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1009
		when "001111110001" => B1 := "1111011"; B2 := "1111110"; B3 := "1111110"; B4 := "0110000"; 
		--1010
		when "001111110010" => B1 := "1111110"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1011
		when "001111110011" => B1 := "0110000"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1012
		when "001111110100" => B1 := "1101101"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1013
		when "001111110101" => B1 := "1111001"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1014
		when "001111110110" => B1 := "0110011"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1015
		when "001111110111" => B1 := "1011011"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1016
		when "001111111000" => B1 := "1011111"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1017
		when "001111111001" => B1 := "1110000"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1018
		when "001111111010" => B1 := "1111111"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1019
		when "001111111011" => B1 := "1111011"; B2 := "0110000"; B3 := "1111110"; B4 := "0110000"; 
		--1020
		when "001111111100" => B1 := "1111110"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1021
		when "001111111101" => B1 := "0110000"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1022
		when "001111111110" => B1 := "1101101"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1023
		when "001111111111" => B1 := "1111001"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1024
		when "010000000000" => B1 := "0110011"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1025
		when "010000000001" => B1 := "1011011"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1026
		when "010000000010" => B1 := "1011111"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1027
		when "010000000011" => B1 := "1110000"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1028
		when "010000000100" => B1 := "1111111"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1029
		when "010000000101" => B1 := "1111011"; B2 := "1101101"; B3 := "1111110"; B4 := "0110000"; 
		--1030
		when "010000000110" => B1 := "1111110"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1031
		when "010000000111" => B1 := "0110000"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1032
		when "010000001000" => B1 := "1101101"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1033
		when "010000001001" => B1 := "1111001"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1034
		when "010000001010" => B1 := "0110011"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1035
		when "010000001011" => B1 := "1011011"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1036
		when "010000001100" => B1 := "1011111"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1037
		when "010000001101" => B1 := "1110000"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1038
		when "010000001110" => B1 := "1111111"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1039
		when "010000001111" => B1 := "1111011"; B2 := "1111001"; B3 := "1111110"; B4 := "0110000"; 
		--1040
		when "010000010000" => B1 := "1111110"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1041
		when "010000010001" => B1 := "0110000"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1042
		when "010000010010" => B1 := "1101101"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1043
		when "010000010011" => B1 := "1111001"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1044
		when "010000010100" => B1 := "0110011"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1045
		when "010000010101" => B1 := "1011011"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1046
		when "010000010110" => B1 := "1011111"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1047
		when "010000010111" => B1 := "1110000"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1048
		when "010000011000" => B1 := "1111111"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1049
		when "010000011001" => B1 := "1111011"; B2 := "0110011"; B3 := "1111110"; B4 := "0110000"; 
		--1050
		when "010000011010" => B1 := "1111110"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1051
		when "010000011011" => B1 := "0110000"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1052
		when "010000011100" => B1 := "1101101"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1053
		when "010000011101" => B1 := "1111001"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1054
		when "010000011110" => B1 := "0110011"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1055
		when "010000011111" => B1 := "1011011"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1056
		when "010000100000" => B1 := "1011111"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1057
		when "010000100001" => B1 := "1110000"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1058
		when "010000100010" => B1 := "1111111"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1059
		when "010000100011" => B1 := "1111011"; B2 := "1011011"; B3 := "1111110"; B4 := "0110000"; 
		--1060
		when "010000100100" => B1 := "1111110"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1061
		when "010000100101" => B1 := "0110000"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1062
		when "010000100110" => B1 := "1101101"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1063
		when "010000100111" => B1 := "1111001"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1064
		when "010000101000" => B1 := "0110011"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1065
		when "010000101001" => B1 := "1011011"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1066
		when "010000101010" => B1 := "1011111"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1067
		when "010000101011" => B1 := "1110000"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1068
		when "010000101100" => B1 := "1111111"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1069
		when "010000101101" => B1 := "1111011"; B2 := "1011111"; B3 := "1111110"; B4 := "0110000"; 
		--1070
		when "010000101110" => B1 := "1111110"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1071
		when "010000101111" => B1 := "0110000"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1072
		when "010000110000" => B1 := "1101101"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1073
		when "010000110001" => B1 := "1111001"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1074
		when "010000110010" => B1 := "0110011"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1075
		when "010000110011" => B1 := "1011011"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1076
		when "010000110100" => B1 := "1011111"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1077
		when "010000110101" => B1 := "1110000"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1078
		when "010000110110" => B1 := "1111111"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1079
		when "010000110111" => B1 := "1111011"; B2 := "1110000"; B3 := "1111110"; B4 := "0110000"; 
		--1080
		when "010000111000" => B1 := "1111110"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1081
		when "010000111001" => B1 := "0110000"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1082
		when "010000111010" => B1 := "1101101"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1083
		when "010000111011" => B1 := "1111001"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1084
		when "010000111100" => B1 := "0110011"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1085
		when "010000111101" => B1 := "1011011"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1086
		when "010000111110" => B1 := "1011111"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1087
		when "010000111111" => B1 := "1110000"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1088
		when "010001000000" => B1 := "1111111"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1089
		when "010001000001" => B1 := "1111011"; B2 := "1111111"; B3 := "1111110"; B4 := "0110000"; 
		--1090
		when "010001000010" => B1 := "1111110"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1091
		when "010001000011" => B1 := "0110000"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1092
		when "010001000100" => B1 := "1101101"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1093
		when "010001000101" => B1 := "1111001"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1094
		when "010001000110" => B1 := "0110011"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1095
		when "010001000111" => B1 := "1011011"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1096
		when "010001001000" => B1 := "1011111"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1097
		when "010001001001" => B1 := "1110000"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1098
		when "010001001010" => B1 := "1111111"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1099
		when "010001001011" => B1 := "1111011"; B2 := "1111011"; B3 := "1111110"; B4 := "0110000"; 
		--1100
		when "010001001100" => B1 := "1111110"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1101
		when "010001001101" => B1 := "0110000"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1102
		when "010001001110" => B1 := "1101101"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1103
		when "010001001111" => B1 := "1111001"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1104
		when "010001010000" => B1 := "0110011"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1105
		when "010001010001" => B1 := "1011011"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1106
		when "010001010010" => B1 := "1011111"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1107
		when "010001010011" => B1 := "1110000"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1108
		when "010001010100" => B1 := "1111111"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1109
		when "010001010101" => B1 := "1111011"; B2 := "1111110"; B3 := "0110000"; B4 := "0110000"; 
		--1110
		when "010001010110" => B1 := "1111110"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1111
		when "010001010111" => B1 := "0110000"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1112
		when "010001011000" => B1 := "1101101"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1113
		when "010001011001" => B1 := "1111001"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1114
		when "010001011010" => B1 := "0110011"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1115
		when "010001011011" => B1 := "1011011"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1116
		when "010001011100" => B1 := "1011111"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1117
		when "010001011101" => B1 := "1110000"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1118
		when "010001011110" => B1 := "1111111"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1119
		when "010001011111" => B1 := "1111011"; B2 := "0110000"; B3 := "0110000"; B4 := "0110000"; 
		--1120
		when "010001100000" => B1 := "1111110"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1121
		when "010001100001" => B1 := "0110000"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1122
		when "010001100010" => B1 := "1101101"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1123
		when "010001100011" => B1 := "1111001"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1124
		when "010001100100" => B1 := "0110011"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1125
		when "010001100101" => B1 := "1011011"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1126
		when "010001100110" => B1 := "1011111"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1127
		when "010001100111" => B1 := "1110000"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1128
		when "010001101000" => B1 := "1111111"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1129
		when "010001101001" => B1 := "1111011"; B2 := "1101101"; B3 := "0110000"; B4 := "0110000"; 
		--1130
		when "010001101010" => B1 := "1111110"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1131
		when "010001101011" => B1 := "0110000"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1132
		when "010001101100" => B1 := "1101101"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1133
		when "010001101101" => B1 := "1111001"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1134
		when "010001101110" => B1 := "0110011"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1135
		when "010001101111" => B1 := "1011011"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1136
		when "010001110000" => B1 := "1011111"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1137
		when "010001110001" => B1 := "1110000"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1138
		when "010001110010" => B1 := "1111111"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1139
		when "010001110011" => B1 := "1111011"; B2 := "1111001"; B3 := "0110000"; B4 := "0110000"; 
		--1140
		when "010001110100" => B1 := "1111110"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1141
		when "010001110101" => B1 := "0110000"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1142
		when "010001110110" => B1 := "1101101"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1143
		when "010001110111" => B1 := "1111001"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1144
		when "010001111000" => B1 := "0110011"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1145
		when "010001111001" => B1 := "1011011"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1146
		when "010001111010" => B1 := "1011111"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1147
		when "010001111011" => B1 := "1110000"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1148
		when "010001111100" => B1 := "1111111"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1149
		when "010001111101" => B1 := "1111011"; B2 := "0110011"; B3 := "0110000"; B4 := "0110000"; 
		--1150
		when "010001111110" => B1 := "1111110"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1151
		when "010001111111" => B1 := "0110000"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1152
		when "010010000000" => B1 := "1101101"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1153
		when "010010000001" => B1 := "1111001"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1154
		when "010010000010" => B1 := "0110011"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1155
		when "010010000011" => B1 := "1011011"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1156
		when "010010000100" => B1 := "1011111"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1157
		when "010010000101" => B1 := "1110000"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1158
		when "010010000110" => B1 := "1111111"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1159
		when "010010000111" => B1 := "1111011"; B2 := "1011011"; B3 := "0110000"; B4 := "0110000"; 
		--1160
		when "010010001000" => B1 := "1111110"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1161
		when "010010001001" => B1 := "0110000"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1162
		when "010010001010" => B1 := "1101101"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1163
		when "010010001011" => B1 := "1111001"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1164
		when "010010001100" => B1 := "0110011"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1165
		when "010010001101" => B1 := "1011011"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1166
		when "010010001110" => B1 := "1011111"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1167
		when "010010001111" => B1 := "1110000"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1168
		when "010010010000" => B1 := "1111111"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1169
		when "010010010001" => B1 := "1111011"; B2 := "1011111"; B3 := "0110000"; B4 := "0110000"; 
		--1170
		when "010010010010" => B1 := "1111110"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1171
		when "010010010011" => B1 := "0110000"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1172
		when "010010010100" => B1 := "1101101"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1173
		when "010010010101" => B1 := "1111001"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1174
		when "010010010110" => B1 := "0110011"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1175
		when "010010010111" => B1 := "1011011"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1176
		when "010010011000" => B1 := "1011111"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1177
		when "010010011001" => B1 := "1110000"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1178
		when "010010011010" => B1 := "1111111"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1179
		when "010010011011" => B1 := "1111011"; B2 := "1110000"; B3 := "0110000"; B4 := "0110000"; 
		--1180
		when "010010011100" => B1 := "1111110"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1181
		when "010010011101" => B1 := "0110000"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1182
		when "010010011110" => B1 := "1101101"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1183
		when "010010011111" => B1 := "1111001"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1184
		when "010010100000" => B1 := "0110011"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1185
		when "010010100001" => B1 := "1011011"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1186
		when "010010100010" => B1 := "1011111"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1187
		when "010010100011" => B1 := "1110000"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1188
		when "010010100100" => B1 := "1111111"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1189
		when "010010100101" => B1 := "1111011"; B2 := "1111111"; B3 := "0110000"; B4 := "0110000"; 
		--1190
		when "010010100110" => B1 := "1111110"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1191
		when "010010100111" => B1 := "0110000"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1192
		when "010010101000" => B1 := "1101101"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1193
		when "010010101001" => B1 := "1111001"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1194
		when "010010101010" => B1 := "0110011"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1195
		when "010010101011" => B1 := "1011011"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1196
		when "010010101100" => B1 := "1011111"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1197
		when "010010101101" => B1 := "1110000"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1198
		when "010010101110" => B1 := "1111111"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1199
		when "010010101111" => B1 := "1111011"; B2 := "1111011"; B3 := "0110000"; B4 := "0110000"; 
		--1200
		when "010010110000" => B1 := "1111110"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1201
		when "010010110001" => B1 := "0110000"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1202
		when "010010110010" => B1 := "1101101"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1203
		when "010010110011" => B1 := "1111001"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1204
		when "010010110100" => B1 := "0110011"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1205
		when "010010110101" => B1 := "1011011"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1206
		when "010010110110" => B1 := "1011111"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1207
		when "010010110111" => B1 := "1110000"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1208
		when "010010111000" => B1 := "1111111"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1209
		when "010010111001" => B1 := "1111011"; B2 := "1111110"; B3 := "1101101"; B4 := "0110000"; 
		--1210
		when "010010111010" => B1 := "1111110"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1211
		when "010010111011" => B1 := "0110000"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1212
		when "010010111100" => B1 := "1101101"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1213
		when "010010111101" => B1 := "1111001"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1214
		when "010010111110" => B1 := "0110011"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1215
		when "010010111111" => B1 := "1011011"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1216
		when "010011000000" => B1 := "1011111"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1217
		when "010011000001" => B1 := "1110000"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1218
		when "010011000010" => B1 := "1111111"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1219
		when "010011000011" => B1 := "1111011"; B2 := "0110000"; B3 := "1101101"; B4 := "0110000"; 
		--1220
		when "010011000100" => B1 := "1111110"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1221
		when "010011000101" => B1 := "0110000"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1222
		when "010011000110" => B1 := "1101101"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1223
		when "010011000111" => B1 := "1111001"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1224
		when "010011001000" => B1 := "0110011"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1225
		when "010011001001" => B1 := "1011011"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1226
		when "010011001010" => B1 := "1011111"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1227
		when "010011001011" => B1 := "1110000"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1228
		when "010011001100" => B1 := "1111111"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1229
		when "010011001101" => B1 := "1111011"; B2 := "1101101"; B3 := "1101101"; B4 := "0110000"; 
		--1230
		when "010011001110" => B1 := "1111110"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1231
		when "010011001111" => B1 := "0110000"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1232
		when "010011010000" => B1 := "1101101"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1233
		when "010011010001" => B1 := "1111001"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1234
		when "010011010010" => B1 := "0110011"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1235
		when "010011010011" => B1 := "1011011"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1236
		when "010011010100" => B1 := "1011111"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1237
		when "010011010101" => B1 := "1110000"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1238
		when "010011010110" => B1 := "1111111"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1239
		when "010011010111" => B1 := "1111011"; B2 := "1111001"; B3 := "1101101"; B4 := "0110000"; 
		--1240
		when "010011011000" => B1 := "1111110"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1241
		when "010011011001" => B1 := "0110000"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1242
		when "010011011010" => B1 := "1101101"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1243
		when "010011011011" => B1 := "1111001"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1244
		when "010011011100" => B1 := "0110011"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1245
		when "010011011101" => B1 := "1011011"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1246
		when "010011011110" => B1 := "1011111"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1247
		when "010011011111" => B1 := "1110000"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1248
		when "010011100000" => B1 := "1111111"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1249
		when "010011100001" => B1 := "1111011"; B2 := "0110011"; B3 := "1101101"; B4 := "0110000"; 
		--1250
		when "010011100010" => B1 := "1111110"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1251
		when "010011100011" => B1 := "0110000"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1252
		when "010011100100" => B1 := "1101101"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1253
		when "010011100101" => B1 := "1111001"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1254
		when "010011100110" => B1 := "0110011"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1255
		when "010011100111" => B1 := "1011011"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1256
		when "010011101000" => B1 := "1011111"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1257
		when "010011101001" => B1 := "1110000"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1258
		when "010011101010" => B1 := "1111111"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1259
		when "010011101011" => B1 := "1111011"; B2 := "1011011"; B3 := "1101101"; B4 := "0110000"; 
		--1260
		when "010011101100" => B1 := "1111110"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1261
		when "010011101101" => B1 := "0110000"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1262
		when "010011101110" => B1 := "1101101"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1263
		when "010011101111" => B1 := "1111001"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1264
		when "010011110000" => B1 := "0110011"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1265
		when "010011110001" => B1 := "1011011"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1266
		when "010011110010" => B1 := "1011111"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1267
		when "010011110011" => B1 := "1110000"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1268
		when "010011110100" => B1 := "1111111"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1269
		when "010011110101" => B1 := "1111011"; B2 := "1011111"; B3 := "1101101"; B4 := "0110000"; 
		--1270
		when "010011110110" => B1 := "1111110"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1271
		when "010011110111" => B1 := "0110000"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1272
		when "010011111000" => B1 := "1101101"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1273
		when "010011111001" => B1 := "1111001"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1274
		when "010011111010" => B1 := "0110011"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1275
		when "010011111011" => B1 := "1011011"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1276
		when "010011111100" => B1 := "1011111"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1277
		when "010011111101" => B1 := "1110000"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1278
		when "010011111110" => B1 := "1111111"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1279
		when "010011111111" => B1 := "1111011"; B2 := "1110000"; B3 := "1101101"; B4 := "0110000"; 
		--1280
		when "010100000000" => B1 := "1111110"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1281
		when "010100000001" => B1 := "0110000"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1282
		when "010100000010" => B1 := "1101101"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1283
		when "010100000011" => B1 := "1111001"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1284
		when "010100000100" => B1 := "0110011"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1285
		when "010100000101" => B1 := "1011011"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1286
		when "010100000110" => B1 := "1011111"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1287
		when "010100000111" => B1 := "1110000"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1288
		when "010100001000" => B1 := "1111111"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1289
		when "010100001001" => B1 := "1111011"; B2 := "1111111"; B3 := "1101101"; B4 := "0110000"; 
		--1290
		when "010100001010" => B1 := "1111110"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1291
		when "010100001011" => B1 := "0110000"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1292
		when "010100001100" => B1 := "1101101"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1293
		when "010100001101" => B1 := "1111001"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1294
		when "010100001110" => B1 := "0110011"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1295
		when "010100001111" => B1 := "1011011"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1296
		when "010100010000" => B1 := "1011111"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1297
		when "010100010001" => B1 := "1110000"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1298
		when "010100010010" => B1 := "1111111"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1299
		when "010100010011" => B1 := "1111011"; B2 := "1111011"; B3 := "1101101"; B4 := "0110000"; 
		--1300
		when "010100010100" => B1 := "1111110"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1301
		when "010100010101" => B1 := "0110000"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1302
		when "010100010110" => B1 := "1101101"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1303
		when "010100010111" => B1 := "1111001"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1304
		when "010100011000" => B1 := "0110011"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1305
		when "010100011001" => B1 := "1011011"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1306
		when "010100011010" => B1 := "1011111"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1307
		when "010100011011" => B1 := "1110000"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1308
		when "010100011100" => B1 := "1111111"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1309
		when "010100011101" => B1 := "1111011"; B2 := "1111110"; B3 := "1111001"; B4 := "0110000"; 
		--1310
		when "010100011110" => B1 := "1111110"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1311
		when "010100011111" => B1 := "0110000"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1312
		when "010100100000" => B1 := "1101101"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1313
		when "010100100001" => B1 := "1111001"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1314
		when "010100100010" => B1 := "0110011"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1315
		when "010100100011" => B1 := "1011011"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1316
		when "010100100100" => B1 := "1011111"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1317
		when "010100100101" => B1 := "1110000"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1318
		when "010100100110" => B1 := "1111111"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1319
		when "010100100111" => B1 := "1111011"; B2 := "0110000"; B3 := "1111001"; B4 := "0110000"; 
		--1320
		when "010100101000" => B1 := "1111110"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1321
		when "010100101001" => B1 := "0110000"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1322
		when "010100101010" => B1 := "1101101"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1323
		when "010100101011" => B1 := "1111001"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1324
		when "010100101100" => B1 := "0110011"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1325
		when "010100101101" => B1 := "1011011"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1326
		when "010100101110" => B1 := "1011111"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1327
		when "010100101111" => B1 := "1110000"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1328
		when "010100110000" => B1 := "1111111"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1329
		when "010100110001" => B1 := "1111011"; B2 := "1101101"; B3 := "1111001"; B4 := "0110000"; 
		--1330
		when "010100110010" => B1 := "1111110"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1331
		when "010100110011" => B1 := "0110000"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1332
		when "010100110100" => B1 := "1101101"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1333
		when "010100110101" => B1 := "1111001"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1334
		when "010100110110" => B1 := "0110011"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1335
		when "010100110111" => B1 := "1011011"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1336
		when "010100111000" => B1 := "1011111"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1337
		when "010100111001" => B1 := "1110000"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1338
		when "010100111010" => B1 := "1111111"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1339
		when "010100111011" => B1 := "1111011"; B2 := "1111001"; B3 := "1111001"; B4 := "0110000"; 
		--1340
		when "010100111100" => B1 := "1111110"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1341
		when "010100111101" => B1 := "0110000"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1342
		when "010100111110" => B1 := "1101101"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1343
		when "010100111111" => B1 := "1111001"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1344
		when "010101000000" => B1 := "0110011"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1345
		when "010101000001" => B1 := "1011011"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1346
		when "010101000010" => B1 := "1011111"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1347
		when "010101000011" => B1 := "1110000"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1348
		when "010101000100" => B1 := "1111111"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1349
		when "010101000101" => B1 := "1111011"; B2 := "0110011"; B3 := "1111001"; B4 := "0110000"; 
		--1350
		when "010101000110" => B1 := "1111110"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1351
		when "010101000111" => B1 := "0110000"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1352
		when "010101001000" => B1 := "1101101"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1353
		when "010101001001" => B1 := "1111001"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1354
		when "010101001010" => B1 := "0110011"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1355
		when "010101001011" => B1 := "1011011"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1356
		when "010101001100" => B1 := "1011111"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1357
		when "010101001101" => B1 := "1110000"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1358
		when "010101001110" => B1 := "1111111"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1359
		when "010101001111" => B1 := "1111011"; B2 := "1011011"; B3 := "1111001"; B4 := "0110000"; 
		--1360
		when "010101010000" => B1 := "1111110"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1361
		when "010101010001" => B1 := "0110000"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1362
		when "010101010010" => B1 := "1101101"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1363
		when "010101010011" => B1 := "1111001"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1364
		when "010101010100" => B1 := "0110011"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1365
		when "010101010101" => B1 := "1011011"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1366
		when "010101010110" => B1 := "1011111"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1367
		when "010101010111" => B1 := "1110000"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1368
		when "010101011000" => B1 := "1111111"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1369
		when "010101011001" => B1 := "1111011"; B2 := "1011111"; B3 := "1111001"; B4 := "0110000"; 
		--1370
		when "010101011010" => B1 := "1111110"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1371
		when "010101011011" => B1 := "0110000"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1372
		when "010101011100" => B1 := "1101101"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1373
		when "010101011101" => B1 := "1111001"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1374
		when "010101011110" => B1 := "0110011"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1375
		when "010101011111" => B1 := "1011011"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1376
		when "010101100000" => B1 := "1011111"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1377
		when "010101100001" => B1 := "1110000"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1378
		when "010101100010" => B1 := "1111111"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1379
		when "010101100011" => B1 := "1111011"; B2 := "1110000"; B3 := "1111001"; B4 := "0110000"; 
		--1380
		when "010101100100" => B1 := "1111110"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1381
		when "010101100101" => B1 := "0110000"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1382
		when "010101100110" => B1 := "1101101"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1383
		when "010101100111" => B1 := "1111001"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1384
		when "010101101000" => B1 := "0110011"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1385
		when "010101101001" => B1 := "1011011"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1386
		when "010101101010" => B1 := "1011111"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1387
		when "010101101011" => B1 := "1110000"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1388
		when "010101101100" => B1 := "1111111"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1389
		when "010101101101" => B1 := "1111011"; B2 := "1111111"; B3 := "1111001"; B4 := "0110000"; 
		--1390
		when "010101101110" => B1 := "1111110"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1391
		when "010101101111" => B1 := "0110000"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1392
		when "010101110000" => B1 := "1101101"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1393
		when "010101110001" => B1 := "1111001"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1394
		when "010101110010" => B1 := "0110011"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1395
		when "010101110011" => B1 := "1011011"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1396
		when "010101110100" => B1 := "1011111"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1397
		when "010101110101" => B1 := "1110000"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1398
		when "010101110110" => B1 := "1111111"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1399
		when "010101110111" => B1 := "1111011"; B2 := "1111011"; B3 := "1111001"; B4 := "0110000"; 
		--1400
		when "010101111000" => B1 := "1111110"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1401
		when "010101111001" => B1 := "0110000"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1402
		when "010101111010" => B1 := "1101101"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1403
		when "010101111011" => B1 := "1111001"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1404
		when "010101111100" => B1 := "0110011"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1405
		when "010101111101" => B1 := "1011011"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1406
		when "010101111110" => B1 := "1011111"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1407
		when "010101111111" => B1 := "1110000"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1408
		when "010110000000" => B1 := "1111111"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1409
		when "010110000001" => B1 := "1111011"; B2 := "1111110"; B3 := "0110011"; B4 := "0110000"; 
		--1410
		when "010110000010" => B1 := "1111110"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1411
		when "010110000011" => B1 := "0110000"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1412
		when "010110000100" => B1 := "1101101"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1413
		when "010110000101" => B1 := "1111001"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1414
		when "010110000110" => B1 := "0110011"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1415
		when "010110000111" => B1 := "1011011"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1416
		when "010110001000" => B1 := "1011111"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1417
		when "010110001001" => B1 := "1110000"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1418
		when "010110001010" => B1 := "1111111"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1419
		when "010110001011" => B1 := "1111011"; B2 := "0110000"; B3 := "0110011"; B4 := "0110000"; 
		--1420
		when "010110001100" => B1 := "1111110"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1421
		when "010110001101" => B1 := "0110000"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1422
		when "010110001110" => B1 := "1101101"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1423
		when "010110001111" => B1 := "1111001"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1424
		when "010110010000" => B1 := "0110011"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1425
		when "010110010001" => B1 := "1011011"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1426
		when "010110010010" => B1 := "1011111"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1427
		when "010110010011" => B1 := "1110000"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1428
		when "010110010100" => B1 := "1111111"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1429
		when "010110010101" => B1 := "1111011"; B2 := "1101101"; B3 := "0110011"; B4 := "0110000"; 
		--1430
		when "010110010110" => B1 := "1111110"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1431
		when "010110010111" => B1 := "0110000"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1432
		when "010110011000" => B1 := "1101101"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1433
		when "010110011001" => B1 := "1111001"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1434
		when "010110011010" => B1 := "0110011"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1435
		when "010110011011" => B1 := "1011011"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1436
		when "010110011100" => B1 := "1011111"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1437
		when "010110011101" => B1 := "1110000"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1438
		when "010110011110" => B1 := "1111111"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1439
		when "010110011111" => B1 := "1111011"; B2 := "1111001"; B3 := "0110011"; B4 := "0110000"; 
		--1440
		when "010110100000" => B1 := "1111110"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1441
		when "010110100001" => B1 := "0110000"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1442
		when "010110100010" => B1 := "1101101"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1443
		when "010110100011" => B1 := "1111001"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1444
		when "010110100100" => B1 := "0110011"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1445
		when "010110100101" => B1 := "1011011"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1446
		when "010110100110" => B1 := "1011111"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1447
		when "010110100111" => B1 := "1110000"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1448
		when "010110101000" => B1 := "1111111"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1449
		when "010110101001" => B1 := "1111011"; B2 := "0110011"; B3 := "0110011"; B4 := "0110000"; 
		--1450
		when "010110101010" => B1 := "1111110"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1451
		when "010110101011" => B1 := "0110000"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1452
		when "010110101100" => B1 := "1101101"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1453
		when "010110101101" => B1 := "1111001"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1454
		when "010110101110" => B1 := "0110011"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1455
		when "010110101111" => B1 := "1011011"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1456
		when "010110110000" => B1 := "1011111"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1457
		when "010110110001" => B1 := "1110000"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1458
		when "010110110010" => B1 := "1111111"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1459
		when "010110110011" => B1 := "1111011"; B2 := "1011011"; B3 := "0110011"; B4 := "0110000"; 
		--1460
		when "010110110100" => B1 := "1111110"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1461
		when "010110110101" => B1 := "0110000"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1462
		when "010110110110" => B1 := "1101101"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1463
		when "010110110111" => B1 := "1111001"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1464
		when "010110111000" => B1 := "0110011"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1465
		when "010110111001" => B1 := "1011011"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1466
		when "010110111010" => B1 := "1011111"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1467
		when "010110111011" => B1 := "1110000"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1468
		when "010110111100" => B1 := "1111111"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1469
		when "010110111101" => B1 := "1111011"; B2 := "1011111"; B3 := "0110011"; B4 := "0110000"; 
		--1470
		when "010110111110" => B1 := "1111110"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1471
		when "010110111111" => B1 := "0110000"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1472
		when "010111000000" => B1 := "1101101"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1473
		when "010111000001" => B1 := "1111001"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1474
		when "010111000010" => B1 := "0110011"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1475
		when "010111000011" => B1 := "1011011"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1476
		when "010111000100" => B1 := "1011111"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1477
		when "010111000101" => B1 := "1110000"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1478
		when "010111000110" => B1 := "1111111"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1479
		when "010111000111" => B1 := "1111011"; B2 := "1110000"; B3 := "0110011"; B4 := "0110000"; 
		--1480
		when "010111001000" => B1 := "1111110"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1481
		when "010111001001" => B1 := "0110000"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1482
		when "010111001010" => B1 := "1101101"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1483
		when "010111001011" => B1 := "1111001"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1484
		when "010111001100" => B1 := "0110011"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1485
		when "010111001101" => B1 := "1011011"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1486
		when "010111001110" => B1 := "1011111"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1487
		when "010111001111" => B1 := "1110000"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1488
		when "010111010000" => B1 := "1111111"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1489
		when "010111010001" => B1 := "1111011"; B2 := "1111111"; B3 := "0110011"; B4 := "0110000"; 
		--1490
		when "010111010010" => B1 := "1111110"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1491
		when "010111010011" => B1 := "0110000"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1492
		when "010111010100" => B1 := "1101101"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1493
		when "010111010101" => B1 := "1111001"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1494
		when "010111010110" => B1 := "0110011"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1495
		when "010111010111" => B1 := "1011011"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1496
		when "010111011000" => B1 := "1011111"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1497
		when "010111011001" => B1 := "1110000"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1498
		when "010111011010" => B1 := "1111111"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1499
		when "010111011011" => B1 := "1111011"; B2 := "1111011"; B3 := "0110011"; B4 := "0110000"; 
		--1500
		when "010111011100" => B1 := "1111110"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1501
		when "010111011101" => B1 := "0110000"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1502
		when "010111011110" => B1 := "1101101"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1503
		when "010111011111" => B1 := "1111001"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1504
		when "010111100000" => B1 := "0110011"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1505
		when "010111100001" => B1 := "1011011"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1506
		when "010111100010" => B1 := "1011111"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1507
		when "010111100011" => B1 := "1110000"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1508
		when "010111100100" => B1 := "1111111"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1509
		when "010111100101" => B1 := "1111011"; B2 := "1111110"; B3 := "1011011"; B4 := "0110000"; 
		--1510
		when "010111100110" => B1 := "1111110"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1511
		when "010111100111" => B1 := "0110000"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1512
		when "010111101000" => B1 := "1101101"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1513
		when "010111101001" => B1 := "1111001"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1514
		when "010111101010" => B1 := "0110011"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1515
		when "010111101011" => B1 := "1011011"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1516
		when "010111101100" => B1 := "1011111"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1517
		when "010111101101" => B1 := "1110000"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1518
		when "010111101110" => B1 := "1111111"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1519
		when "010111101111" => B1 := "1111011"; B2 := "0110000"; B3 := "1011011"; B4 := "0110000"; 
		--1520
		when "010111110000" => B1 := "1111110"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1521
		when "010111110001" => B1 := "0110000"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1522
		when "010111110010" => B1 := "1101101"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1523
		when "010111110011" => B1 := "1111001"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1524
		when "010111110100" => B1 := "0110011"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1525
		when "010111110101" => B1 := "1011011"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1526
		when "010111110110" => B1 := "1011111"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1527
		when "010111110111" => B1 := "1110000"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1528
		when "010111111000" => B1 := "1111111"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1529
		when "010111111001" => B1 := "1111011"; B2 := "1101101"; B3 := "1011011"; B4 := "0110000"; 
		--1530
		when "010111111010" => B1 := "1111110"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1531
		when "010111111011" => B1 := "0110000"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1532
		when "010111111100" => B1 := "1101101"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1533
		when "010111111101" => B1 := "1111001"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1534
		when "010111111110" => B1 := "0110011"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1535
		when "010111111111" => B1 := "1011011"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1536
		when "011000000000" => B1 := "1011111"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1537
		when "011000000001" => B1 := "1110000"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1538
		when "011000000010" => B1 := "1111111"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1539
		when "011000000011" => B1 := "1111011"; B2 := "1111001"; B3 := "1011011"; B4 := "0110000"; 
		--1540
		when "011000000100" => B1 := "1111110"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1541
		when "011000000101" => B1 := "0110000"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1542
		when "011000000110" => B1 := "1101101"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1543
		when "011000000111" => B1 := "1111001"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1544
		when "011000001000" => B1 := "0110011"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1545
		when "011000001001" => B1 := "1011011"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1546
		when "011000001010" => B1 := "1011111"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1547
		when "011000001011" => B1 := "1110000"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1548
		when "011000001100" => B1 := "1111111"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1549
		when "011000001101" => B1 := "1111011"; B2 := "0110011"; B3 := "1011011"; B4 := "0110000"; 
		--1550
		when "011000001110" => B1 := "1111110"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1551
		when "011000001111" => B1 := "0110000"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1552
		when "011000010000" => B1 := "1101101"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1553
		when "011000010001" => B1 := "1111001"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1554
		when "011000010010" => B1 := "0110011"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1555
		when "011000010011" => B1 := "1011011"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1556
		when "011000010100" => B1 := "1011111"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1557
		when "011000010101" => B1 := "1110000"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1558
		when "011000010110" => B1 := "1111111"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1559
		when "011000010111" => B1 := "1111011"; B2 := "1011011"; B3 := "1011011"; B4 := "0110000"; 
		--1560
		when "011000011000" => B1 := "1111110"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1561
		when "011000011001" => B1 := "0110000"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1562
		when "011000011010" => B1 := "1101101"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1563
		when "011000011011" => B1 := "1111001"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1564
		when "011000011100" => B1 := "0110011"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1565
		when "011000011101" => B1 := "1011011"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1566
		when "011000011110" => B1 := "1011111"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1567
		when "011000011111" => B1 := "1110000"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1568
		when "011000100000" => B1 := "1111111"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1569
		when "011000100001" => B1 := "1111011"; B2 := "1011111"; B3 := "1011011"; B4 := "0110000"; 
		--1570
		when "011000100010" => B1 := "1111110"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1571
		when "011000100011" => B1 := "0110000"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1572
		when "011000100100" => B1 := "1101101"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1573
		when "011000100101" => B1 := "1111001"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1574
		when "011000100110" => B1 := "0110011"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1575
		when "011000100111" => B1 := "1011011"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1576
		when "011000101000" => B1 := "1011111"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1577
		when "011000101001" => B1 := "1110000"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1578
		when "011000101010" => B1 := "1111111"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1579
		when "011000101011" => B1 := "1111011"; B2 := "1110000"; B3 := "1011011"; B4 := "0110000"; 
		--1580
		when "011000101100" => B1 := "1111110"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1581
		when "011000101101" => B1 := "0110000"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1582
		when "011000101110" => B1 := "1101101"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1583
		when "011000101111" => B1 := "1111001"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1584
		when "011000110000" => B1 := "0110011"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1585
		when "011000110001" => B1 := "1011011"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1586
		when "011000110010" => B1 := "1011111"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1587
		when "011000110011" => B1 := "1110000"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1588
		when "011000110100" => B1 := "1111111"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1589
		when "011000110101" => B1 := "1111011"; B2 := "1111111"; B3 := "1011011"; B4 := "0110000"; 
		--1590
		when "011000110110" => B1 := "1111110"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1591
		when "011000110111" => B1 := "0110000"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1592
		when "011000111000" => B1 := "1101101"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1593
		when "011000111001" => B1 := "1111001"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1594
		when "011000111010" => B1 := "0110011"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1595
		when "011000111011" => B1 := "1011011"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1596
		when "011000111100" => B1 := "1011111"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1597
		when "011000111101" => B1 := "1110000"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1598
		when "011000111110" => B1 := "1111111"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1599
		when "011000111111" => B1 := "1111011"; B2 := "1111011"; B3 := "1011011"; B4 := "0110000"; 
		--1600
		when "011001000000" => B1 := "1111110"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1601
		when "011001000001" => B1 := "0110000"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1602
		when "011001000010" => B1 := "1101101"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1603
		when "011001000011" => B1 := "1111001"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1604
		when "011001000100" => B1 := "0110011"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1605
		when "011001000101" => B1 := "1011011"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1606
		when "011001000110" => B1 := "1011111"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1607
		when "011001000111" => B1 := "1110000"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1608
		when "011001001000" => B1 := "1111111"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1609
		when "011001001001" => B1 := "1111011"; B2 := "1111110"; B3 := "1011111"; B4 := "0110000"; 
		--1610
		when "011001001010" => B1 := "1111110"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1611
		when "011001001011" => B1 := "0110000"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1612
		when "011001001100" => B1 := "1101101"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1613
		when "011001001101" => B1 := "1111001"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1614
		when "011001001110" => B1 := "0110011"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1615
		when "011001001111" => B1 := "1011011"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1616
		when "011001010000" => B1 := "1011111"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1617
		when "011001010001" => B1 := "1110000"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1618
		when "011001010010" => B1 := "1111111"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1619
		when "011001010011" => B1 := "1111011"; B2 := "0110000"; B3 := "1011111"; B4 := "0110000"; 
		--1620
		when "011001010100" => B1 := "1111110"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1621
		when "011001010101" => B1 := "0110000"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1622
		when "011001010110" => B1 := "1101101"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1623
		when "011001010111" => B1 := "1111001"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1624
		when "011001011000" => B1 := "0110011"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1625
		when "011001011001" => B1 := "1011011"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1626
		when "011001011010" => B1 := "1011111"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1627
		when "011001011011" => B1 := "1110000"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1628
		when "011001011100" => B1 := "1111111"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1629
		when "011001011101" => B1 := "1111011"; B2 := "1101101"; B3 := "1011111"; B4 := "0110000"; 
		--1630
		when "011001011110" => B1 := "1111110"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1631
		when "011001011111" => B1 := "0110000"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1632
		when "011001100000" => B1 := "1101101"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1633
		when "011001100001" => B1 := "1111001"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1634
		when "011001100010" => B1 := "0110011"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1635
		when "011001100011" => B1 := "1011011"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1636
		when "011001100100" => B1 := "1011111"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1637
		when "011001100101" => B1 := "1110000"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1638
		when "011001100110" => B1 := "1111111"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1639
		when "011001100111" => B1 := "1111011"; B2 := "1111001"; B3 := "1011111"; B4 := "0110000"; 
		--1640
		when "011001101000" => B1 := "1111110"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1641
		when "011001101001" => B1 := "0110000"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1642
		when "011001101010" => B1 := "1101101"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1643
		when "011001101011" => B1 := "1111001"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1644
		when "011001101100" => B1 := "0110011"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1645
		when "011001101101" => B1 := "1011011"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1646
		when "011001101110" => B1 := "1011111"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1647
		when "011001101111" => B1 := "1110000"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1648
		when "011001110000" => B1 := "1111111"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1649
		when "011001110001" => B1 := "1111011"; B2 := "0110011"; B3 := "1011111"; B4 := "0110000"; 
		--1650
		when "011001110010" => B1 := "1111110"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1651
		when "011001110011" => B1 := "0110000"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1652
		when "011001110100" => B1 := "1101101"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1653
		when "011001110101" => B1 := "1111001"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1654
		when "011001110110" => B1 := "0110011"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1655
		when "011001110111" => B1 := "1011011"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1656
		when "011001111000" => B1 := "1011111"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1657
		when "011001111001" => B1 := "1110000"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1658
		when "011001111010" => B1 := "1111111"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1659
		when "011001111011" => B1 := "1111011"; B2 := "1011011"; B3 := "1011111"; B4 := "0110000"; 
		--1660
		when "011001111100" => B1 := "1111110"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1661
		when "011001111101" => B1 := "0110000"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1662
		when "011001111110" => B1 := "1101101"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1663
		when "011001111111" => B1 := "1111001"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1664
		when "011010000000" => B1 := "0110011"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1665
		when "011010000001" => B1 := "1011011"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1666
		when "011010000010" => B1 := "1011111"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1667
		when "011010000011" => B1 := "1110000"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1668
		when "011010000100" => B1 := "1111111"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1669
		when "011010000101" => B1 := "1111011"; B2 := "1011111"; B3 := "1011111"; B4 := "0110000"; 
		--1670
		when "011010000110" => B1 := "1111110"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1671
		when "011010000111" => B1 := "0110000"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1672
		when "011010001000" => B1 := "1101101"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1673
		when "011010001001" => B1 := "1111001"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1674
		when "011010001010" => B1 := "0110011"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1675
		when "011010001011" => B1 := "1011011"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1676
		when "011010001100" => B1 := "1011111"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1677
		when "011010001101" => B1 := "1110000"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1678
		when "011010001110" => B1 := "1111111"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1679
		when "011010001111" => B1 := "1111011"; B2 := "1110000"; B3 := "1011111"; B4 := "0110000"; 
		--1680
		when "011010010000" => B1 := "1111110"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1681
		when "011010010001" => B1 := "0110000"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1682
		when "011010010010" => B1 := "1101101"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1683
		when "011010010011" => B1 := "1111001"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1684
		when "011010010100" => B1 := "0110011"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1685
		when "011010010101" => B1 := "1011011"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1686
		when "011010010110" => B1 := "1011111"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1687
		when "011010010111" => B1 := "1110000"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1688
		when "011010011000" => B1 := "1111111"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1689
		when "011010011001" => B1 := "1111011"; B2 := "1111111"; B3 := "1011111"; B4 := "0110000"; 
		--1690
		when "011010011010" => B1 := "1111110"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1691
		when "011010011011" => B1 := "0110000"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1692
		when "011010011100" => B1 := "1101101"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1693
		when "011010011101" => B1 := "1111001"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1694
		when "011010011110" => B1 := "0110011"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1695
		when "011010011111" => B1 := "1011011"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1696
		when "011010100000" => B1 := "1011111"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1697
		when "011010100001" => B1 := "1110000"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1698
		when "011010100010" => B1 := "1111111"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1699
		when "011010100011" => B1 := "1111011"; B2 := "1111011"; B3 := "1011111"; B4 := "0110000"; 
		--1700
		when "011010100100" => B1 := "1111110"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1701
		when "011010100101" => B1 := "0110000"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1702
		when "011010100110" => B1 := "1101101"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1703
		when "011010100111" => B1 := "1111001"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1704
		when "011010101000" => B1 := "0110011"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1705
		when "011010101001" => B1 := "1011011"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1706
		when "011010101010" => B1 := "1011111"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1707
		when "011010101011" => B1 := "1110000"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1708
		when "011010101100" => B1 := "1111111"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1709
		when "011010101101" => B1 := "1111011"; B2 := "1111110"; B3 := "1110000"; B4 := "0110000"; 
		--1710
		when "011010101110" => B1 := "1111110"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1711
		when "011010101111" => B1 := "0110000"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1712
		when "011010110000" => B1 := "1101101"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1713
		when "011010110001" => B1 := "1111001"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1714
		when "011010110010" => B1 := "0110011"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1715
		when "011010110011" => B1 := "1011011"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1716
		when "011010110100" => B1 := "1011111"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1717
		when "011010110101" => B1 := "1110000"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1718
		when "011010110110" => B1 := "1111111"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1719
		when "011010110111" => B1 := "1111011"; B2 := "0110000"; B3 := "1110000"; B4 := "0110000"; 
		--1720
		when "011010111000" => B1 := "1111110"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1721
		when "011010111001" => B1 := "0110000"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1722
		when "011010111010" => B1 := "1101101"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1723
		when "011010111011" => B1 := "1111001"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1724
		when "011010111100" => B1 := "0110011"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1725
		when "011010111101" => B1 := "1011011"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1726
		when "011010111110" => B1 := "1011111"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1727
		when "011010111111" => B1 := "1110000"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1728
		when "011011000000" => B1 := "1111111"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1729
		when "011011000001" => B1 := "1111011"; B2 := "1101101"; B3 := "1110000"; B4 := "0110000"; 
		--1730
		when "011011000010" => B1 := "1111110"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1731
		when "011011000011" => B1 := "0110000"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1732
		when "011011000100" => B1 := "1101101"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1733
		when "011011000101" => B1 := "1111001"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1734
		when "011011000110" => B1 := "0110011"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1735
		when "011011000111" => B1 := "1011011"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1736
		when "011011001000" => B1 := "1011111"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1737
		when "011011001001" => B1 := "1110000"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1738
		when "011011001010" => B1 := "1111111"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1739
		when "011011001011" => B1 := "1111011"; B2 := "1111001"; B3 := "1110000"; B4 := "0110000"; 
		--1740
		when "011011001100" => B1 := "1111110"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1741
		when "011011001101" => B1 := "0110000"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1742
		when "011011001110" => B1 := "1101101"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1743
		when "011011001111" => B1 := "1111001"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1744
		when "011011010000" => B1 := "0110011"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1745
		when "011011010001" => B1 := "1011011"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1746
		when "011011010010" => B1 := "1011111"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1747
		when "011011010011" => B1 := "1110000"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1748
		when "011011010100" => B1 := "1111111"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1749
		when "011011010101" => B1 := "1111011"; B2 := "0110011"; B3 := "1110000"; B4 := "0110000"; 
		--1750
		when "011011010110" => B1 := "1111110"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1751
		when "011011010111" => B1 := "0110000"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1752
		when "011011011000" => B1 := "1101101"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1753
		when "011011011001" => B1 := "1111001"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1754
		when "011011011010" => B1 := "0110011"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1755
		when "011011011011" => B1 := "1011011"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1756
		when "011011011100" => B1 := "1011111"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1757
		when "011011011101" => B1 := "1110000"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1758
		when "011011011110" => B1 := "1111111"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1759
		when "011011011111" => B1 := "1111011"; B2 := "1011011"; B3 := "1110000"; B4 := "0110000"; 
		--1760
		when "011011100000" => B1 := "1111110"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1761
		when "011011100001" => B1 := "0110000"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1762
		when "011011100010" => B1 := "1101101"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1763
		when "011011100011" => B1 := "1111001"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1764
		when "011011100100" => B1 := "0110011"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1765
		when "011011100101" => B1 := "1011011"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1766
		when "011011100110" => B1 := "1011111"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1767
		when "011011100111" => B1 := "1110000"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1768
		when "011011101000" => B1 := "1111111"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1769
		when "011011101001" => B1 := "1111011"; B2 := "1011111"; B3 := "1110000"; B4 := "0110000"; 
		--1770
		when "011011101010" => B1 := "1111110"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1771
		when "011011101011" => B1 := "0110000"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1772
		when "011011101100" => B1 := "1101101"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1773
		when "011011101101" => B1 := "1111001"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1774
		when "011011101110" => B1 := "0110011"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1775
		when "011011101111" => B1 := "1011011"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1776
		when "011011110000" => B1 := "1011111"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1777
		when "011011110001" => B1 := "1110000"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1778
		when "011011110010" => B1 := "1111111"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1779
		when "011011110011" => B1 := "1111011"; B2 := "1110000"; B3 := "1110000"; B4 := "0110000"; 
		--1780
		when "011011110100" => B1 := "1111110"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1781
		when "011011110101" => B1 := "0110000"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1782
		when "011011110110" => B1 := "1101101"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1783
		when "011011110111" => B1 := "1111001"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1784
		when "011011111000" => B1 := "0110011"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1785
		when "011011111001" => B1 := "1011011"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1786
		when "011011111010" => B1 := "1011111"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1787
		when "011011111011" => B1 := "1110000"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1788
		when "011011111100" => B1 := "1111111"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1789
		when "011011111101" => B1 := "1111011"; B2 := "1111111"; B3 := "1110000"; B4 := "0110000"; 
		--1790
		when "011011111110" => B1 := "1111110"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1791
		when "011011111111" => B1 := "0110000"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1792
		when "011100000000" => B1 := "1101101"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1793
		when "011100000001" => B1 := "1111001"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1794
		when "011100000010" => B1 := "0110011"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1795
		when "011100000011" => B1 := "1011011"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1796
		when "011100000100" => B1 := "1011111"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1797
		when "011100000101" => B1 := "1110000"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1798
		when "011100000110" => B1 := "1111111"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1799
		when "011100000111" => B1 := "1111011"; B2 := "1111011"; B3 := "1110000"; B4 := "0110000"; 
		--1800
		when "011100001000" => B1 := "1111110"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1801
		when "011100001001" => B1 := "0110000"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1802
		when "011100001010" => B1 := "1101101"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1803
		when "011100001011" => B1 := "1111001"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1804
		when "011100001100" => B1 := "0110011"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1805
		when "011100001101" => B1 := "1011011"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1806
		when "011100001110" => B1 := "1011111"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1807
		when "011100001111" => B1 := "1110000"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1808
		when "011100010000" => B1 := "1111111"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1809
		when "011100010001" => B1 := "1111011"; B2 := "1111110"; B3 := "1111111"; B4 := "0110000"; 
		--1810
		when "011100010010" => B1 := "1111110"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1811
		when "011100010011" => B1 := "0110000"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1812
		when "011100010100" => B1 := "1101101"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1813
		when "011100010101" => B1 := "1111001"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1814
		when "011100010110" => B1 := "0110011"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1815
		when "011100010111" => B1 := "1011011"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1816
		when "011100011000" => B1 := "1011111"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1817
		when "011100011001" => B1 := "1110000"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1818
		when "011100011010" => B1 := "1111111"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1819
		when "011100011011" => B1 := "1111011"; B2 := "0110000"; B3 := "1111111"; B4 := "0110000"; 
		--1820
		when "011100011100" => B1 := "1111110"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1821
		when "011100011101" => B1 := "0110000"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1822
		when "011100011110" => B1 := "1101101"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1823
		when "011100011111" => B1 := "1111001"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1824
		when "011100100000" => B1 := "0110011"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1825
		when "011100100001" => B1 := "1011011"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1826
		when "011100100010" => B1 := "1011111"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1827
		when "011100100011" => B1 := "1110000"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1828
		when "011100100100" => B1 := "1111111"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1829
		when "011100100101" => B1 := "1111011"; B2 := "1101101"; B3 := "1111111"; B4 := "0110000"; 
		--1830
		when "011100100110" => B1 := "1111110"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1831
		when "011100100111" => B1 := "0110000"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1832
		when "011100101000" => B1 := "1101101"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1833
		when "011100101001" => B1 := "1111001"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1834
		when "011100101010" => B1 := "0110011"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1835
		when "011100101011" => B1 := "1011011"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1836
		when "011100101100" => B1 := "1011111"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1837
		when "011100101101" => B1 := "1110000"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1838
		when "011100101110" => B1 := "1111111"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1839
		when "011100101111" => B1 := "1111011"; B2 := "1111001"; B3 := "1111111"; B4 := "0110000"; 
		--1840
		when "011100110000" => B1 := "1111110"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1841
		when "011100110001" => B1 := "0110000"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1842
		when "011100110010" => B1 := "1101101"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1843
		when "011100110011" => B1 := "1111001"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1844
		when "011100110100" => B1 := "0110011"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1845
		when "011100110101" => B1 := "1011011"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1846
		when "011100110110" => B1 := "1011111"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1847
		when "011100110111" => B1 := "1110000"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1848
		when "011100111000" => B1 := "1111111"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1849
		when "011100111001" => B1 := "1111011"; B2 := "0110011"; B3 := "1111111"; B4 := "0110000"; 
		--1850
		when "011100111010" => B1 := "1111110"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1851
		when "011100111011" => B1 := "0110000"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1852
		when "011100111100" => B1 := "1101101"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1853
		when "011100111101" => B1 := "1111001"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1854
		when "011100111110" => B1 := "0110011"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1855
		when "011100111111" => B1 := "1011011"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1856
		when "011101000000" => B1 := "1011111"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1857
		when "011101000001" => B1 := "1110000"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1858
		when "011101000010" => B1 := "1111111"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1859
		when "011101000011" => B1 := "1111011"; B2 := "1011011"; B3 := "1111111"; B4 := "0110000"; 
		--1860
		when "011101000100" => B1 := "1111110"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1861
		when "011101000101" => B1 := "0110000"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1862
		when "011101000110" => B1 := "1101101"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1863
		when "011101000111" => B1 := "1111001"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1864
		when "011101001000" => B1 := "0110011"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1865
		when "011101001001" => B1 := "1011011"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1866
		when "011101001010" => B1 := "1011111"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1867
		when "011101001011" => B1 := "1110000"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1868
		when "011101001100" => B1 := "1111111"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1869
		when "011101001101" => B1 := "1111011"; B2 := "1011111"; B3 := "1111111"; B4 := "0110000"; 
		--1870
		when "011101001110" => B1 := "1111110"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1871
		when "011101001111" => B1 := "0110000"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1872
		when "011101010000" => B1 := "1101101"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1873
		when "011101010001" => B1 := "1111001"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1874
		when "011101010010" => B1 := "0110011"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1875
		when "011101010011" => B1 := "1011011"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1876
		when "011101010100" => B1 := "1011111"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1877
		when "011101010101" => B1 := "1110000"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1878
		when "011101010110" => B1 := "1111111"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1879
		when "011101010111" => B1 := "1111011"; B2 := "1110000"; B3 := "1111111"; B4 := "0110000"; 
		--1880
		when "011101011000" => B1 := "1111110"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1881
		when "011101011001" => B1 := "0110000"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1882
		when "011101011010" => B1 := "1101101"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1883
		when "011101011011" => B1 := "1111001"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1884
		when "011101011100" => B1 := "0110011"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1885
		when "011101011101" => B1 := "1011011"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1886
		when "011101011110" => B1 := "1011111"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1887
		when "011101011111" => B1 := "1110000"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1888
		when "011101100000" => B1 := "1111111"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1889
		when "011101100001" => B1 := "1111011"; B2 := "1111111"; B3 := "1111111"; B4 := "0110000"; 
		--1890
		when "011101100010" => B1 := "1111110"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1891
		when "011101100011" => B1 := "0110000"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1892
		when "011101100100" => B1 := "1101101"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1893
		when "011101100101" => B1 := "1111001"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1894
		when "011101100110" => B1 := "0110011"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1895
		when "011101100111" => B1 := "1011011"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1896
		when "011101101000" => B1 := "1011111"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1897
		when "011101101001" => B1 := "1110000"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1898
		when "011101101010" => B1 := "1111111"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1899
		when "011101101011" => B1 := "1111011"; B2 := "1111011"; B3 := "1111111"; B4 := "0110000"; 
		--1900
		when "011101101100" => B1 := "1111110"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1901
		when "011101101101" => B1 := "0110000"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1902
		when "011101101110" => B1 := "1101101"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1903
		when "011101101111" => B1 := "1111001"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1904
		when "011101110000" => B1 := "0110011"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1905
		when "011101110001" => B1 := "1011011"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1906
		when "011101110010" => B1 := "1011111"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1907
		when "011101110011" => B1 := "1110000"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1908
		when "011101110100" => B1 := "1111111"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1909
		when "011101110101" => B1 := "1111011"; B2 := "1111110"; B3 := "1111011"; B4 := "0110000"; 
		--1910
		when "011101110110" => B1 := "1111110"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1911
		when "011101110111" => B1 := "0110000"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1912
		when "011101111000" => B1 := "1101101"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1913
		when "011101111001" => B1 := "1111001"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1914
		when "011101111010" => B1 := "0110011"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1915
		when "011101111011" => B1 := "1011011"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1916
		when "011101111100" => B1 := "1011111"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1917
		when "011101111101" => B1 := "1110000"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1918
		when "011101111110" => B1 := "1111111"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1919
		when "011101111111" => B1 := "1111011"; B2 := "0110000"; B3 := "1111011"; B4 := "0110000"; 
		--1920
		when "011110000000" => B1 := "1111110"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1921
		when "011110000001" => B1 := "0110000"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1922
		when "011110000010" => B1 := "1101101"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1923
		when "011110000011" => B1 := "1111001"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1924
		when "011110000100" => B1 := "0110011"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1925
		when "011110000101" => B1 := "1011011"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1926
		when "011110000110" => B1 := "1011111"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1927
		when "011110000111" => B1 := "1110000"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1928
		when "011110001000" => B1 := "1111111"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1929
		when "011110001001" => B1 := "1111011"; B2 := "1101101"; B3 := "1111011"; B4 := "0110000"; 
		--1930
		when "011110001010" => B1 := "1111110"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1931
		when "011110001011" => B1 := "0110000"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1932
		when "011110001100" => B1 := "1101101"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1933
		when "011110001101" => B1 := "1111001"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1934
		when "011110001110" => B1 := "0110011"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1935
		when "011110001111" => B1 := "1011011"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1936
		when "011110010000" => B1 := "1011111"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1937
		when "011110010001" => B1 := "1110000"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1938
		when "011110010010" => B1 := "1111111"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1939
		when "011110010011" => B1 := "1111011"; B2 := "1111001"; B3 := "1111011"; B4 := "0110000"; 
		--1940
		when "011110010100" => B1 := "1111110"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1941
		when "011110010101" => B1 := "0110000"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1942
		when "011110010110" => B1 := "1101101"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1943
		when "011110010111" => B1 := "1111001"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1944
		when "011110011000" => B1 := "0110011"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1945
		when "011110011001" => B1 := "1011011"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1946
		when "011110011010" => B1 := "1011111"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1947
		when "011110011011" => B1 := "1110000"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1948
		when "011110011100" => B1 := "1111111"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1949
		when "011110011101" => B1 := "1111011"; B2 := "0110011"; B3 := "1111011"; B4 := "0110000"; 
		--1950
		when "011110011110" => B1 := "1111110"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1951
		when "011110011111" => B1 := "0110000"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1952
		when "011110100000" => B1 := "1101101"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1953
		when "011110100001" => B1 := "1111001"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1954
		when "011110100010" => B1 := "0110011"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1955
		when "011110100011" => B1 := "1011011"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1956
		when "011110100100" => B1 := "1011111"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1957
		when "011110100101" => B1 := "1110000"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1958
		when "011110100110" => B1 := "1111111"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1959
		when "011110100111" => B1 := "1111011"; B2 := "1011011"; B3 := "1111011"; B4 := "0110000"; 
		--1960
		when "011110101000" => B1 := "1111110"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1961
		when "011110101001" => B1 := "0110000"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1962
		when "011110101010" => B1 := "1101101"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1963
		when "011110101011" => B1 := "1111001"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1964
		when "011110101100" => B1 := "0110011"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1965
		when "011110101101" => B1 := "1011011"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1966
		when "011110101110" => B1 := "1011111"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1967
		when "011110101111" => B1 := "1110000"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1968
		when "011110110000" => B1 := "1111111"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1969
		when "011110110001" => B1 := "1111011"; B2 := "1011111"; B3 := "1111011"; B4 := "0110000"; 
		--1970
		when "011110110010" => B1 := "1111110"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1971
		when "011110110011" => B1 := "0110000"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1972
		when "011110110100" => B1 := "1101101"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1973
		when "011110110101" => B1 := "1111001"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1974
		when "011110110110" => B1 := "0110011"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1975
		when "011110110111" => B1 := "1011011"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1976
		when "011110111000" => B1 := "1011111"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1977
		when "011110111001" => B1 := "1110000"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1978
		when "011110111010" => B1 := "1111111"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1979
		when "011110111011" => B1 := "1111011"; B2 := "1110000"; B3 := "1111011"; B4 := "0110000"; 
		--1980
		when "011110111100" => B1 := "1111110"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1981
		when "011110111101" => B1 := "0110000"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1982
		when "011110111110" => B1 := "1101101"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1983
		when "011110111111" => B1 := "1111001"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1984
		when "011111000000" => B1 := "0110011"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1985
		when "011111000001" => B1 := "1011011"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1986
		when "011111000010" => B1 := "1011111"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1987
		when "011111000011" => B1 := "1110000"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1988
		when "011111000100" => B1 := "1111111"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1989
		when "011111000101" => B1 := "1111011"; B2 := "1111111"; B3 := "1111011"; B4 := "0110000"; 
		--1990
		when "011111000110" => B1 := "1111110"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--1991
		when "011111000111" => B1 := "0110000"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--1992
		when "011111001000" => B1 := "1101101"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--1993
		when "011111001001" => B1 := "1111001"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--1994
		when "011111001010" => B1 := "0110011"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--1995
		when "011111001011" => B1 := "1011011"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--1996
		when "011111001100" => B1 := "1011111"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--1997
		when "011111001101" => B1 := "1110000"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--1998
		when "011111001110" => B1 := "1111111"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--1999
		when "011111001111" => B1 := "1111011"; B2 := "1111011"; B3 := "1111011"; B4 := "0110000"; 
		--2000
		when "011111010000" => B1 := "1111110"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2001
		when "011111010001" => B1 := "0110000"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2002
		when "011111010010" => B1 := "1101101"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2003
		when "011111010011" => B1 := "1111001"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2004
		when "011111010100" => B1 := "0110011"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2005
		when "011111010101" => B1 := "1011011"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2006
		when "011111010110" => B1 := "1011111"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2007
		when "011111010111" => B1 := "1110000"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2008
		when "011111011000" => B1 := "1111111"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2009
		when "011111011001" => B1 := "1111011"; B2 := "1111110"; B3 := "1111110"; B4 := "1101101"; 
		--2010
		when "011111011010" => B1 := "1111110"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2011
		when "011111011011" => B1 := "0110000"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2012
		when "011111011100" => B1 := "1101101"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2013
		when "011111011101" => B1 := "1111001"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2014
		when "011111011110" => B1 := "0110011"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2015
		when "011111011111" => B1 := "1011011"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2016
		when "011111100000" => B1 := "1011111"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2017
		when "011111100001" => B1 := "1110000"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2018
		when "011111100010" => B1 := "1111111"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2019
		when "011111100011" => B1 := "1111011"; B2 := "0110000"; B3 := "1111110"; B4 := "1101101"; 
		--2020
		when "011111100100" => B1 := "1111110"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2021
		when "011111100101" => B1 := "0110000"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2022
		when "011111100110" => B1 := "1101101"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2023
		when "011111100111" => B1 := "1111001"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2024
		when "011111101000" => B1 := "0110011"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2025
		when "011111101001" => B1 := "1011011"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2026
		when "011111101010" => B1 := "1011111"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2027
		when "011111101011" => B1 := "1110000"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2028
		when "011111101100" => B1 := "1111111"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2029
		when "011111101101" => B1 := "1111011"; B2 := "1101101"; B3 := "1111110"; B4 := "1101101"; 
		--2030
		when "011111101110" => B1 := "1111110"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2031
		when "011111101111" => B1 := "0110000"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2032
		when "011111110000" => B1 := "1101101"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2033
		when "011111110001" => B1 := "1111001"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2034
		when "011111110010" => B1 := "0110011"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2035
		when "011111110011" => B1 := "1011011"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2036
		when "011111110100" => B1 := "1011111"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2037
		when "011111110101" => B1 := "1110000"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2038
		when "011111110110" => B1 := "1111111"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2039
		when "011111110111" => B1 := "1111011"; B2 := "1111001"; B3 := "1111110"; B4 := "1101101"; 
		--2040
		when "011111111000" => B1 := "1111110"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2041
		when "011111111001" => B1 := "0110000"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2042
		when "011111111010" => B1 := "1101101"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2043
		when "011111111011" => B1 := "1111001"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2044
		when "011111111100" => B1 := "0110011"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2045
		when "011111111101" => B1 := "1011011"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2046
		when "011111111110" => B1 := "1011111"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2047
		when "011111111111" => B1 := "1110000"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2048
		when "100000000000" => B1 := "1111111"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2049
		when "100000000001" => B1 := "1111011"; B2 := "0110011"; B3 := "1111110"; B4 := "1101101"; 
		--2050
		when "100000000010" => B1 := "1111110"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2051
		when "100000000011" => B1 := "0110000"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2052
		when "100000000100" => B1 := "1101101"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2053
		when "100000000101" => B1 := "1111001"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2054
		when "100000000110" => B1 := "0110011"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2055
		when "100000000111" => B1 := "1011011"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2056
		when "100000001000" => B1 := "1011111"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2057
		when "100000001001" => B1 := "1110000"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2058
		when "100000001010" => B1 := "1111111"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2059
		when "100000001011" => B1 := "1111011"; B2 := "1011011"; B3 := "1111110"; B4 := "1101101"; 
		--2060
		when "100000001100" => B1 := "1111110"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2061
		when "100000001101" => B1 := "0110000"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2062
		when "100000001110" => B1 := "1101101"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2063
		when "100000001111" => B1 := "1111001"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2064
		when "100000010000" => B1 := "0110011"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2065
		when "100000010001" => B1 := "1011011"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2066
		when "100000010010" => B1 := "1011111"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2067
		when "100000010011" => B1 := "1110000"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2068
		when "100000010100" => B1 := "1111111"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2069
		when "100000010101" => B1 := "1111011"; B2 := "1011111"; B3 := "1111110"; B4 := "1101101"; 
		--2070
		when "100000010110" => B1 := "1111110"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2071
		when "100000010111" => B1 := "0110000"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2072
		when "100000011000" => B1 := "1101101"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2073
		when "100000011001" => B1 := "1111001"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2074
		when "100000011010" => B1 := "0110011"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2075
		when "100000011011" => B1 := "1011011"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2076
		when "100000011100" => B1 := "1011111"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2077
		when "100000011101" => B1 := "1110000"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2078
		when "100000011110" => B1 := "1111111"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2079
		when "100000011111" => B1 := "1111011"; B2 := "1110000"; B3 := "1111110"; B4 := "1101101"; 
		--2080
		when "100000100000" => B1 := "1111110"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2081
		when "100000100001" => B1 := "0110000"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2082
		when "100000100010" => B1 := "1101101"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2083
		when "100000100011" => B1 := "1111001"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2084
		when "100000100100" => B1 := "0110011"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2085
		when "100000100101" => B1 := "1011011"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2086
		when "100000100110" => B1 := "1011111"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2087
		when "100000100111" => B1 := "1110000"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2088
		when "100000101000" => B1 := "1111111"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2089
		when "100000101001" => B1 := "1111011"; B2 := "1111111"; B3 := "1111110"; B4 := "1101101"; 
		--2090
		when "100000101010" => B1 := "1111110"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2091
		when "100000101011" => B1 := "0110000"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2092
		when "100000101100" => B1 := "1101101"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2093
		when "100000101101" => B1 := "1111001"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2094
		when "100000101110" => B1 := "0110011"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2095
		when "100000101111" => B1 := "1011011"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2096
		when "100000110000" => B1 := "1011111"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2097
		when "100000110001" => B1 := "1110000"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2098
		when "100000110010" => B1 := "1111111"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2099
		when "100000110011" => B1 := "1111011"; B2 := "1111011"; B3 := "1111110"; B4 := "1101101"; 
		--2100
		when "100000110100" => B1 := "1111110"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2101
		when "100000110101" => B1 := "0110000"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2102
		when "100000110110" => B1 := "1101101"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2103
		when "100000110111" => B1 := "1111001"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2104
		when "100000111000" => B1 := "0110011"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2105
		when "100000111001" => B1 := "1011011"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2106
		when "100000111010" => B1 := "1011111"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2107
		when "100000111011" => B1 := "1110000"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2108
		when "100000111100" => B1 := "1111111"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2109
		when "100000111101" => B1 := "1111011"; B2 := "1111110"; B3 := "0110000"; B4 := "1101101"; 
		--2110
		when "100000111110" => B1 := "1111110"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2111
		when "100000111111" => B1 := "0110000"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2112
		when "100001000000" => B1 := "1101101"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2113
		when "100001000001" => B1 := "1111001"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2114
		when "100001000010" => B1 := "0110011"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2115
		when "100001000011" => B1 := "1011011"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2116
		when "100001000100" => B1 := "1011111"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2117
		when "100001000101" => B1 := "1110000"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2118
		when "100001000110" => B1 := "1111111"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2119
		when "100001000111" => B1 := "1111011"; B2 := "0110000"; B3 := "0110000"; B4 := "1101101"; 
		--2120
		when "100001001000" => B1 := "1111110"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2121
		when "100001001001" => B1 := "0110000"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2122
		when "100001001010" => B1 := "1101101"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2123
		when "100001001011" => B1 := "1111001"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2124
		when "100001001100" => B1 := "0110011"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2125
		when "100001001101" => B1 := "1011011"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2126
		when "100001001110" => B1 := "1011111"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2127
		when "100001001111" => B1 := "1110000"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2128
		when "100001010000" => B1 := "1111111"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2129
		when "100001010001" => B1 := "1111011"; B2 := "1101101"; B3 := "0110000"; B4 := "1101101"; 
		--2130
		when "100001010010" => B1 := "1111110"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2131
		when "100001010011" => B1 := "0110000"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2132
		when "100001010100" => B1 := "1101101"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2133
		when "100001010101" => B1 := "1111001"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2134
		when "100001010110" => B1 := "0110011"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2135
		when "100001010111" => B1 := "1011011"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2136
		when "100001011000" => B1 := "1011111"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2137
		when "100001011001" => B1 := "1110000"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2138
		when "100001011010" => B1 := "1111111"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2139
		when "100001011011" => B1 := "1111011"; B2 := "1111001"; B3 := "0110000"; B4 := "1101101"; 
		--2140
		when "100001011100" => B1 := "1111110"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2141
		when "100001011101" => B1 := "0110000"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2142
		when "100001011110" => B1 := "1101101"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2143
		when "100001011111" => B1 := "1111001"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2144
		when "100001100000" => B1 := "0110011"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2145
		when "100001100001" => B1 := "1011011"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2146
		when "100001100010" => B1 := "1011111"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2147
		when "100001100011" => B1 := "1110000"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2148
		when "100001100100" => B1 := "1111111"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2149
		when "100001100101" => B1 := "1111011"; B2 := "0110011"; B3 := "0110000"; B4 := "1101101"; 
		--2150
		when "100001100110" => B1 := "1111110"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2151
		when "100001100111" => B1 := "0110000"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2152
		when "100001101000" => B1 := "1101101"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2153
		when "100001101001" => B1 := "1111001"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2154
		when "100001101010" => B1 := "0110011"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2155
		when "100001101011" => B1 := "1011011"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2156
		when "100001101100" => B1 := "1011111"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2157
		when "100001101101" => B1 := "1110000"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2158
		when "100001101110" => B1 := "1111111"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2159
		when "100001101111" => B1 := "1111011"; B2 := "1011011"; B3 := "0110000"; B4 := "1101101"; 
		--2160
		when "100001110000" => B1 := "1111110"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2161
		when "100001110001" => B1 := "0110000"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2162
		when "100001110010" => B1 := "1101101"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2163
		when "100001110011" => B1 := "1111001"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2164
		when "100001110100" => B1 := "0110011"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2165
		when "100001110101" => B1 := "1011011"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2166
		when "100001110110" => B1 := "1011111"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2167
		when "100001110111" => B1 := "1110000"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2168
		when "100001111000" => B1 := "1111111"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2169
		when "100001111001" => B1 := "1111011"; B2 := "1011111"; B3 := "0110000"; B4 := "1101101"; 
		--2170
		when "100001111010" => B1 := "1111110"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2171
		when "100001111011" => B1 := "0110000"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2172
		when "100001111100" => B1 := "1101101"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2173
		when "100001111101" => B1 := "1111001"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2174
		when "100001111110" => B1 := "0110011"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2175
		when "100001111111" => B1 := "1011011"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2176
		when "100010000000" => B1 := "1011111"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2177
		when "100010000001" => B1 := "1110000"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2178
		when "100010000010" => B1 := "1111111"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2179
		when "100010000011" => B1 := "1111011"; B2 := "1110000"; B3 := "0110000"; B4 := "1101101"; 
		--2180
		when "100010000100" => B1 := "1111110"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2181
		when "100010000101" => B1 := "0110000"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2182
		when "100010000110" => B1 := "1101101"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2183
		when "100010000111" => B1 := "1111001"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2184
		when "100010001000" => B1 := "0110011"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2185
		when "100010001001" => B1 := "1011011"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2186
		when "100010001010" => B1 := "1011111"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2187
		when "100010001011" => B1 := "1110000"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2188
		when "100010001100" => B1 := "1111111"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2189
		when "100010001101" => B1 := "1111011"; B2 := "1111111"; B3 := "0110000"; B4 := "1101101"; 
		--2190
		when "100010001110" => B1 := "1111110"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2191
		when "100010001111" => B1 := "0110000"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2192
		when "100010010000" => B1 := "1101101"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2193
		when "100010010001" => B1 := "1111001"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2194
		when "100010010010" => B1 := "0110011"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2195
		when "100010010011" => B1 := "1011011"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2196
		when "100010010100" => B1 := "1011111"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2197
		when "100010010101" => B1 := "1110000"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2198
		when "100010010110" => B1 := "1111111"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2199
		when "100010010111" => B1 := "1111011"; B2 := "1111011"; B3 := "0110000"; B4 := "1101101"; 
		--2200
		when "100010011000" => B1 := "1111110"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2201
		when "100010011001" => B1 := "0110000"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2202
		when "100010011010" => B1 := "1101101"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2203
		when "100010011011" => B1 := "1111001"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2204
		when "100010011100" => B1 := "0110011"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2205
		when "100010011101" => B1 := "1011011"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2206
		when "100010011110" => B1 := "1011111"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2207
		when "100010011111" => B1 := "1110000"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2208
		when "100010100000" => B1 := "1111111"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2209
		when "100010100001" => B1 := "1111011"; B2 := "1111110"; B3 := "1101101"; B4 := "1101101"; 
		--2210
		when "100010100010" => B1 := "1111110"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2211
		when "100010100011" => B1 := "0110000"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2212
		when "100010100100" => B1 := "1101101"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2213
		when "100010100101" => B1 := "1111001"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2214
		when "100010100110" => B1 := "0110011"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2215
		when "100010100111" => B1 := "1011011"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2216
		when "100010101000" => B1 := "1011111"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2217
		when "100010101001" => B1 := "1110000"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2218
		when "100010101010" => B1 := "1111111"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2219
		when "100010101011" => B1 := "1111011"; B2 := "0110000"; B3 := "1101101"; B4 := "1101101"; 
		--2220
		when "100010101100" => B1 := "1111110"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2221
		when "100010101101" => B1 := "0110000"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2222
		when "100010101110" => B1 := "1101101"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2223
		when "100010101111" => B1 := "1111001"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2224
		when "100010110000" => B1 := "0110011"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2225
		when "100010110001" => B1 := "1011011"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2226
		when "100010110010" => B1 := "1011111"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2227
		when "100010110011" => B1 := "1110000"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2228
		when "100010110100" => B1 := "1111111"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2229
		when "100010110101" => B1 := "1111011"; B2 := "1101101"; B3 := "1101101"; B4 := "1101101"; 
		--2230
		when "100010110110" => B1 := "1111110"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2231
		when "100010110111" => B1 := "0110000"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2232
		when "100010111000" => B1 := "1101101"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2233
		when "100010111001" => B1 := "1111001"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2234
		when "100010111010" => B1 := "0110011"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2235
		when "100010111011" => B1 := "1011011"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2236
		when "100010111100" => B1 := "1011111"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2237
		when "100010111101" => B1 := "1110000"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2238
		when "100010111110" => B1 := "1111111"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2239
		when "100010111111" => B1 := "1111011"; B2 := "1111001"; B3 := "1101101"; B4 := "1101101"; 
		--2240
		when "100011000000" => B1 := "1111110"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2241
		when "100011000001" => B1 := "0110000"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2242
		when "100011000010" => B1 := "1101101"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2243
		when "100011000011" => B1 := "1111001"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2244
		when "100011000100" => B1 := "0110011"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2245
		when "100011000101" => B1 := "1011011"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2246
		when "100011000110" => B1 := "1011111"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2247
		when "100011000111" => B1 := "1110000"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2248
		when "100011001000" => B1 := "1111111"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2249
		when "100011001001" => B1 := "1111011"; B2 := "0110011"; B3 := "1101101"; B4 := "1101101"; 
		--2250
		when "100011001010" => B1 := "1111110"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2251
		when "100011001011" => B1 := "0110000"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2252
		when "100011001100" => B1 := "1101101"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2253
		when "100011001101" => B1 := "1111001"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2254
		when "100011001110" => B1 := "0110011"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2255
		when "100011001111" => B1 := "1011011"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2256
		when "100011010000" => B1 := "1011111"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2257
		when "100011010001" => B1 := "1110000"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2258
		when "100011010010" => B1 := "1111111"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2259
		when "100011010011" => B1 := "1111011"; B2 := "1011011"; B3 := "1101101"; B4 := "1101101"; 
		--2260
		when "100011010100" => B1 := "1111110"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2261
		when "100011010101" => B1 := "0110000"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2262
		when "100011010110" => B1 := "1101101"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2263
		when "100011010111" => B1 := "1111001"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2264
		when "100011011000" => B1 := "0110011"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2265
		when "100011011001" => B1 := "1011011"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2266
		when "100011011010" => B1 := "1011111"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2267
		when "100011011011" => B1 := "1110000"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2268
		when "100011011100" => B1 := "1111111"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2269
		when "100011011101" => B1 := "1111011"; B2 := "1011111"; B3 := "1101101"; B4 := "1101101"; 
		--2270
		when "100011011110" => B1 := "1111110"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2271
		when "100011011111" => B1 := "0110000"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2272
		when "100011100000" => B1 := "1101101"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2273
		when "100011100001" => B1 := "1111001"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2274
		when "100011100010" => B1 := "0110011"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2275
		when "100011100011" => B1 := "1011011"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2276
		when "100011100100" => B1 := "1011111"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2277
		when "100011100101" => B1 := "1110000"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2278
		when "100011100110" => B1 := "1111111"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2279
		when "100011100111" => B1 := "1111011"; B2 := "1110000"; B3 := "1101101"; B4 := "1101101"; 
		--2280
		when "100011101000" => B1 := "1111110"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2281
		when "100011101001" => B1 := "0110000"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2282
		when "100011101010" => B1 := "1101101"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2283
		when "100011101011" => B1 := "1111001"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2284
		when "100011101100" => B1 := "0110011"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2285
		when "100011101101" => B1 := "1011011"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2286
		when "100011101110" => B1 := "1011111"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2287
		when "100011101111" => B1 := "1110000"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2288
		when "100011110000" => B1 := "1111111"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2289
		when "100011110001" => B1 := "1111011"; B2 := "1111111"; B3 := "1101101"; B4 := "1101101"; 
		--2290
		when "100011110010" => B1 := "1111110"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2291
		when "100011110011" => B1 := "0110000"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2292
		when "100011110100" => B1 := "1101101"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2293
		when "100011110101" => B1 := "1111001"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2294
		when "100011110110" => B1 := "0110011"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2295
		when "100011110111" => B1 := "1011011"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2296
		when "100011111000" => B1 := "1011111"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2297
		when "100011111001" => B1 := "1110000"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2298
		when "100011111010" => B1 := "1111111"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2299
		when "100011111011" => B1 := "1111011"; B2 := "1111011"; B3 := "1101101"; B4 := "1101101"; 
		--2300
		when "100011111100" => B1 := "1111110"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2301
		when "100011111101" => B1 := "0110000"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2302
		when "100011111110" => B1 := "1101101"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2303
		when "100011111111" => B1 := "1111001"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2304
		when "100100000000" => B1 := "0110011"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2305
		when "100100000001" => B1 := "1011011"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2306
		when "100100000010" => B1 := "1011111"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2307
		when "100100000011" => B1 := "1110000"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2308
		when "100100000100" => B1 := "1111111"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2309
		when "100100000101" => B1 := "1111011"; B2 := "1111110"; B3 := "1111001"; B4 := "1101101"; 
		--2310
		when "100100000110" => B1 := "1111110"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2311
		when "100100000111" => B1 := "0110000"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2312
		when "100100001000" => B1 := "1101101"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2313
		when "100100001001" => B1 := "1111001"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2314
		when "100100001010" => B1 := "0110011"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2315
		when "100100001011" => B1 := "1011011"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2316
		when "100100001100" => B1 := "1011111"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2317
		when "100100001101" => B1 := "1110000"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2318
		when "100100001110" => B1 := "1111111"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2319
		when "100100001111" => B1 := "1111011"; B2 := "0110000"; B3 := "1111001"; B4 := "1101101"; 
		--2320
		when "100100010000" => B1 := "1111110"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2321
		when "100100010001" => B1 := "0110000"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2322
		when "100100010010" => B1 := "1101101"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2323
		when "100100010011" => B1 := "1111001"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2324
		when "100100010100" => B1 := "0110011"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2325
		when "100100010101" => B1 := "1011011"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2326
		when "100100010110" => B1 := "1011111"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2327
		when "100100010111" => B1 := "1110000"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2328
		when "100100011000" => B1 := "1111111"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2329
		when "100100011001" => B1 := "1111011"; B2 := "1101101"; B3 := "1111001"; B4 := "1101101"; 
		--2330
		when "100100011010" => B1 := "1111110"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2331
		when "100100011011" => B1 := "0110000"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2332
		when "100100011100" => B1 := "1101101"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2333
		when "100100011101" => B1 := "1111001"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2334
		when "100100011110" => B1 := "0110011"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2335
		when "100100011111" => B1 := "1011011"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2336
		when "100100100000" => B1 := "1011111"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2337
		when "100100100001" => B1 := "1110000"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2338
		when "100100100010" => B1 := "1111111"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2339
		when "100100100011" => B1 := "1111011"; B2 := "1111001"; B3 := "1111001"; B4 := "1101101"; 
		--2340
		when "100100100100" => B1 := "1111110"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2341
		when "100100100101" => B1 := "0110000"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2342
		when "100100100110" => B1 := "1101101"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2343
		when "100100100111" => B1 := "1111001"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2344
		when "100100101000" => B1 := "0110011"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2345
		when "100100101001" => B1 := "1011011"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2346
		when "100100101010" => B1 := "1011111"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2347
		when "100100101011" => B1 := "1110000"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2348
		when "100100101100" => B1 := "1111111"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2349
		when "100100101101" => B1 := "1111011"; B2 := "0110011"; B3 := "1111001"; B4 := "1101101"; 
		--2350
		when "100100101110" => B1 := "1111110"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2351
		when "100100101111" => B1 := "0110000"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2352
		when "100100110000" => B1 := "1101101"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2353
		when "100100110001" => B1 := "1111001"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2354
		when "100100110010" => B1 := "0110011"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2355
		when "100100110011" => B1 := "1011011"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2356
		when "100100110100" => B1 := "1011111"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2357
		when "100100110101" => B1 := "1110000"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2358
		when "100100110110" => B1 := "1111111"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2359
		when "100100110111" => B1 := "1111011"; B2 := "1011011"; B3 := "1111001"; B4 := "1101101"; 
		--2360
		when "100100111000" => B1 := "1111110"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2361
		when "100100111001" => B1 := "0110000"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2362
		when "100100111010" => B1 := "1101101"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2363
		when "100100111011" => B1 := "1111001"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2364
		when "100100111100" => B1 := "0110011"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2365
		when "100100111101" => B1 := "1011011"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2366
		when "100100111110" => B1 := "1011111"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2367
		when "100100111111" => B1 := "1110000"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2368
		when "100101000000" => B1 := "1111111"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2369
		when "100101000001" => B1 := "1111011"; B2 := "1011111"; B3 := "1111001"; B4 := "1101101"; 
		--2370
		when "100101000010" => B1 := "1111110"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2371
		when "100101000011" => B1 := "0110000"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2372
		when "100101000100" => B1 := "1101101"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2373
		when "100101000101" => B1 := "1111001"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2374
		when "100101000110" => B1 := "0110011"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2375
		when "100101000111" => B1 := "1011011"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2376
		when "100101001000" => B1 := "1011111"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2377
		when "100101001001" => B1 := "1110000"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2378
		when "100101001010" => B1 := "1111111"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2379
		when "100101001011" => B1 := "1111011"; B2 := "1110000"; B3 := "1111001"; B4 := "1101101"; 
		--2380
		when "100101001100" => B1 := "1111110"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2381
		when "100101001101" => B1 := "0110000"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2382
		when "100101001110" => B1 := "1101101"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2383
		when "100101001111" => B1 := "1111001"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2384
		when "100101010000" => B1 := "0110011"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2385
		when "100101010001" => B1 := "1011011"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2386
		when "100101010010" => B1 := "1011111"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2387
		when "100101010011" => B1 := "1110000"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2388
		when "100101010100" => B1 := "1111111"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2389
		when "100101010101" => B1 := "1111011"; B2 := "1111111"; B3 := "1111001"; B4 := "1101101"; 
		--2390
		when "100101010110" => B1 := "1111110"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2391
		when "100101010111" => B1 := "0110000"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2392
		when "100101011000" => B1 := "1101101"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2393
		when "100101011001" => B1 := "1111001"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2394
		when "100101011010" => B1 := "0110011"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2395
		when "100101011011" => B1 := "1011011"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2396
		when "100101011100" => B1 := "1011111"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2397
		when "100101011101" => B1 := "1110000"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2398
		when "100101011110" => B1 := "1111111"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2399
		when "100101011111" => B1 := "1111011"; B2 := "1111011"; B3 := "1111001"; B4 := "1101101"; 
		--2400
		when "100101100000" => B1 := "1111110"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2401
		when "100101100001" => B1 := "0110000"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2402
		when "100101100010" => B1 := "1101101"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2403
		when "100101100011" => B1 := "1111001"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2404
		when "100101100100" => B1 := "0110011"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2405
		when "100101100101" => B1 := "1011011"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2406
		when "100101100110" => B1 := "1011111"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2407
		when "100101100111" => B1 := "1110000"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2408
		when "100101101000" => B1 := "1111111"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2409
		when "100101101001" => B1 := "1111011"; B2 := "1111110"; B3 := "0110011"; B4 := "1101101"; 
		--2410
		when "100101101010" => B1 := "1111110"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2411
		when "100101101011" => B1 := "0110000"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2412
		when "100101101100" => B1 := "1101101"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2413
		when "100101101101" => B1 := "1111001"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2414
		when "100101101110" => B1 := "0110011"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2415
		when "100101101111" => B1 := "1011011"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2416
		when "100101110000" => B1 := "1011111"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2417
		when "100101110001" => B1 := "1110000"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2418
		when "100101110010" => B1 := "1111111"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2419
		when "100101110011" => B1 := "1111011"; B2 := "0110000"; B3 := "0110011"; B4 := "1101101"; 
		--2420
		when "100101110100" => B1 := "1111110"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2421
		when "100101110101" => B1 := "0110000"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2422
		when "100101110110" => B1 := "1101101"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2423
		when "100101110111" => B1 := "1111001"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2424
		when "100101111000" => B1 := "0110011"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2425
		when "100101111001" => B1 := "1011011"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2426
		when "100101111010" => B1 := "1011111"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2427
		when "100101111011" => B1 := "1110000"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2428
		when "100101111100" => B1 := "1111111"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2429
		when "100101111101" => B1 := "1111011"; B2 := "1101101"; B3 := "0110011"; B4 := "1101101"; 
		--2430
		when "100101111110" => B1 := "1111110"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2431
		when "100101111111" => B1 := "0110000"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2432
		when "100110000000" => B1 := "1101101"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2433
		when "100110000001" => B1 := "1111001"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2434
		when "100110000010" => B1 := "0110011"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2435
		when "100110000011" => B1 := "1011011"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2436
		when "100110000100" => B1 := "1011111"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2437
		when "100110000101" => B1 := "1110000"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2438
		when "100110000110" => B1 := "1111111"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2439
		when "100110000111" => B1 := "1111011"; B2 := "1111001"; B3 := "0110011"; B4 := "1101101"; 
		--2440
		when "100110001000" => B1 := "1111110"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2441
		when "100110001001" => B1 := "0110000"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2442
		when "100110001010" => B1 := "1101101"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2443
		when "100110001011" => B1 := "1111001"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2444
		when "100110001100" => B1 := "0110011"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2445
		when "100110001101" => B1 := "1011011"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2446
		when "100110001110" => B1 := "1011111"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2447
		when "100110001111" => B1 := "1110000"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2448
		when "100110010000" => B1 := "1111111"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2449
		when "100110010001" => B1 := "1111011"; B2 := "0110011"; B3 := "0110011"; B4 := "1101101"; 
		--2450
		when "100110010010" => B1 := "1111110"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2451
		when "100110010011" => B1 := "0110000"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2452
		when "100110010100" => B1 := "1101101"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2453
		when "100110010101" => B1 := "1111001"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2454
		when "100110010110" => B1 := "0110011"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2455
		when "100110010111" => B1 := "1011011"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2456
		when "100110011000" => B1 := "1011111"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2457
		when "100110011001" => B1 := "1110000"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2458
		when "100110011010" => B1 := "1111111"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2459
		when "100110011011" => B1 := "1111011"; B2 := "1011011"; B3 := "0110011"; B4 := "1101101"; 
		--2460
		when "100110011100" => B1 := "1111110"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2461
		when "100110011101" => B1 := "0110000"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2462
		when "100110011110" => B1 := "1101101"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2463
		when "100110011111" => B1 := "1111001"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2464
		when "100110100000" => B1 := "0110011"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2465
		when "100110100001" => B1 := "1011011"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2466
		when "100110100010" => B1 := "1011111"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2467
		when "100110100011" => B1 := "1110000"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2468
		when "100110100100" => B1 := "1111111"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2469
		when "100110100101" => B1 := "1111011"; B2 := "1011111"; B3 := "0110011"; B4 := "1101101"; 
		--2470
		when "100110100110" => B1 := "1111110"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2471
		when "100110100111" => B1 := "0110000"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2472
		when "100110101000" => B1 := "1101101"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2473
		when "100110101001" => B1 := "1111001"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2474
		when "100110101010" => B1 := "0110011"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2475
		when "100110101011" => B1 := "1011011"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2476
		when "100110101100" => B1 := "1011111"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2477
		when "100110101101" => B1 := "1110000"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2478
		when "100110101110" => B1 := "1111111"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2479
		when "100110101111" => B1 := "1111011"; B2 := "1110000"; B3 := "0110011"; B4 := "1101101"; 
		--2480
		when "100110110000" => B1 := "1111110"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2481
		when "100110110001" => B1 := "0110000"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2482
		when "100110110010" => B1 := "1101101"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2483
		when "100110110011" => B1 := "1111001"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2484
		when "100110110100" => B1 := "0110011"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2485
		when "100110110101" => B1 := "1011011"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2486
		when "100110110110" => B1 := "1011111"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2487
		when "100110110111" => B1 := "1110000"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2488
		when "100110111000" => B1 := "1111111"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2489
		when "100110111001" => B1 := "1111011"; B2 := "1111111"; B3 := "0110011"; B4 := "1101101"; 
		--2490
		when "100110111010" => B1 := "1111110"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2491
		when "100110111011" => B1 := "0110000"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2492
		when "100110111100" => B1 := "1101101"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2493
		when "100110111101" => B1 := "1111001"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2494
		when "100110111110" => B1 := "0110011"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2495
		when "100110111111" => B1 := "1011011"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2496
		when "100111000000" => B1 := "1011111"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2497
		when "100111000001" => B1 := "1110000"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2498
		when "100111000010" => B1 := "1111111"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2499
		when "100111000011" => B1 := "1111011"; B2 := "1111011"; B3 := "0110011"; B4 := "1101101"; 
		--2500
		when "100111000100" => B1 := "1111110"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2501
		when "100111000101" => B1 := "0110000"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2502
		when "100111000110" => B1 := "1101101"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2503
		when "100111000111" => B1 := "1111001"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2504
		when "100111001000" => B1 := "0110011"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2505
		when "100111001001" => B1 := "1011011"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2506
		when "100111001010" => B1 := "1011111"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2507
		when "100111001011" => B1 := "1110000"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2508
		when "100111001100" => B1 := "1111111"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2509
		when "100111001101" => B1 := "1111011"; B2 := "1111110"; B3 := "1011011"; B4 := "1101101"; 
		--2510
		when "100111001110" => B1 := "1111110"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2511
		when "100111001111" => B1 := "0110000"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2512
		when "100111010000" => B1 := "1101101"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2513
		when "100111010001" => B1 := "1111001"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2514
		when "100111010010" => B1 := "0110011"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2515
		when "100111010011" => B1 := "1011011"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2516
		when "100111010100" => B1 := "1011111"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2517
		when "100111010101" => B1 := "1110000"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2518
		when "100111010110" => B1 := "1111111"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2519
		when "100111010111" => B1 := "1111011"; B2 := "0110000"; B3 := "1011011"; B4 := "1101101"; 
		--2520
		when "100111011000" => B1 := "1111110"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2521
		when "100111011001" => B1 := "0110000"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2522
		when "100111011010" => B1 := "1101101"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2523
		when "100111011011" => B1 := "1111001"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2524
		when "100111011100" => B1 := "0110011"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2525
		when "100111011101" => B1 := "1011011"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2526
		when "100111011110" => B1 := "1011111"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2527
		when "100111011111" => B1 := "1110000"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2528
		when "100111100000" => B1 := "1111111"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2529
		when "100111100001" => B1 := "1111011"; B2 := "1101101"; B3 := "1011011"; B4 := "1101101"; 
		--2530
		when "100111100010" => B1 := "1111110"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2531
		when "100111100011" => B1 := "0110000"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2532
		when "100111100100" => B1 := "1101101"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2533
		when "100111100101" => B1 := "1111001"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2534
		when "100111100110" => B1 := "0110011"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2535
		when "100111100111" => B1 := "1011011"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2536
		when "100111101000" => B1 := "1011111"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2537
		when "100111101001" => B1 := "1110000"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2538
		when "100111101010" => B1 := "1111111"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2539
		when "100111101011" => B1 := "1111011"; B2 := "1111001"; B3 := "1011011"; B4 := "1101101"; 
		--2540
		when "100111101100" => B1 := "1111110"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2541
		when "100111101101" => B1 := "0110000"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2542
		when "100111101110" => B1 := "1101101"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2543
		when "100111101111" => B1 := "1111001"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2544
		when "100111110000" => B1 := "0110011"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2545
		when "100111110001" => B1 := "1011011"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2546
		when "100111110010" => B1 := "1011111"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2547
		when "100111110011" => B1 := "1110000"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2548
		when "100111110100" => B1 := "1111111"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2549
		when "100111110101" => B1 := "1111011"; B2 := "0110011"; B3 := "1011011"; B4 := "1101101"; 
		--2550
		when "100111110110" => B1 := "1111110"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2551
		when "100111110111" => B1 := "0110000"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2552
		when "100111111000" => B1 := "1101101"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2553
		when "100111111001" => B1 := "1111001"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2554
		when "100111111010" => B1 := "0110011"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2555
		when "100111111011" => B1 := "1011011"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2556
		when "100111111100" => B1 := "1011111"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2557
		when "100111111101" => B1 := "1110000"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2558
		when "100111111110" => B1 := "1111111"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2559
		when "100111111111" => B1 := "1111011"; B2 := "1011011"; B3 := "1011011"; B4 := "1101101"; 
		--2560
		when "101000000000" => B1 := "1111110"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2561
		when "101000000001" => B1 := "0110000"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2562
		when "101000000010" => B1 := "1101101"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2563
		when "101000000011" => B1 := "1111001"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2564
		when "101000000100" => B1 := "0110011"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2565
		when "101000000101" => B1 := "1011011"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2566
		when "101000000110" => B1 := "1011111"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2567
		when "101000000111" => B1 := "1110000"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2568
		when "101000001000" => B1 := "1111111"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2569
		when "101000001001" => B1 := "1111011"; B2 := "1011111"; B3 := "1011011"; B4 := "1101101"; 
		--2570
		when "101000001010" => B1 := "1111110"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2571
		when "101000001011" => B1 := "0110000"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2572
		when "101000001100" => B1 := "1101101"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2573
		when "101000001101" => B1 := "1111001"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2574
		when "101000001110" => B1 := "0110011"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2575
		when "101000001111" => B1 := "1011011"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2576
		when "101000010000" => B1 := "1011111"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2577
		when "101000010001" => B1 := "1110000"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2578
		when "101000010010" => B1 := "1111111"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2579
		when "101000010011" => B1 := "1111011"; B2 := "1110000"; B3 := "1011011"; B4 := "1101101"; 
		--2580
		when "101000010100" => B1 := "1111110"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2581
		when "101000010101" => B1 := "0110000"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2582
		when "101000010110" => B1 := "1101101"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2583
		when "101000010111" => B1 := "1111001"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2584
		when "101000011000" => B1 := "0110011"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2585
		when "101000011001" => B1 := "1011011"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2586
		when "101000011010" => B1 := "1011111"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2587
		when "101000011011" => B1 := "1110000"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2588
		when "101000011100" => B1 := "1111111"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2589
		when "101000011101" => B1 := "1111011"; B2 := "1111111"; B3 := "1011011"; B4 := "1101101"; 
		--2590
		when "101000011110" => B1 := "1111110"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2591
		when "101000011111" => B1 := "0110000"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2592
		when "101000100000" => B1 := "1101101"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2593
		when "101000100001" => B1 := "1111001"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2594
		when "101000100010" => B1 := "0110011"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2595
		when "101000100011" => B1 := "1011011"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2596
		when "101000100100" => B1 := "1011111"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2597
		when "101000100101" => B1 := "1110000"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2598
		when "101000100110" => B1 := "1111111"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2599
		when "101000100111" => B1 := "1111011"; B2 := "1111011"; B3 := "1011011"; B4 := "1101101"; 
		--2600
		when "101000101000" => B1 := "1111110"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2601
		when "101000101001" => B1 := "0110000"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2602
		when "101000101010" => B1 := "1101101"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2603
		when "101000101011" => B1 := "1111001"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2604
		when "101000101100" => B1 := "0110011"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2605
		when "101000101101" => B1 := "1011011"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2606
		when "101000101110" => B1 := "1011111"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2607
		when "101000101111" => B1 := "1110000"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2608
		when "101000110000" => B1 := "1111111"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2609
		when "101000110001" => B1 := "1111011"; B2 := "1111110"; B3 := "1011111"; B4 := "1101101"; 
		--2610
		when "101000110010" => B1 := "1111110"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2611
		when "101000110011" => B1 := "0110000"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2612
		when "101000110100" => B1 := "1101101"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2613
		when "101000110101" => B1 := "1111001"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2614
		when "101000110110" => B1 := "0110011"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2615
		when "101000110111" => B1 := "1011011"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2616
		when "101000111000" => B1 := "1011111"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2617
		when "101000111001" => B1 := "1110000"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2618
		when "101000111010" => B1 := "1111111"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2619
		when "101000111011" => B1 := "1111011"; B2 := "0110000"; B3 := "1011111"; B4 := "1101101"; 
		--2620
		when "101000111100" => B1 := "1111110"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2621
		when "101000111101" => B1 := "0110000"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2622
		when "101000111110" => B1 := "1101101"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2623
		when "101000111111" => B1 := "1111001"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2624
		when "101001000000" => B1 := "0110011"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2625
		when "101001000001" => B1 := "1011011"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2626
		when "101001000010" => B1 := "1011111"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2627
		when "101001000011" => B1 := "1110000"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2628
		when "101001000100" => B1 := "1111111"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2629
		when "101001000101" => B1 := "1111011"; B2 := "1101101"; B3 := "1011111"; B4 := "1101101"; 
		--2630
		when "101001000110" => B1 := "1111110"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2631
		when "101001000111" => B1 := "0110000"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2632
		when "101001001000" => B1 := "1101101"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2633
		when "101001001001" => B1 := "1111001"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2634
		when "101001001010" => B1 := "0110011"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2635
		when "101001001011" => B1 := "1011011"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2636
		when "101001001100" => B1 := "1011111"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2637
		when "101001001101" => B1 := "1110000"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2638
		when "101001001110" => B1 := "1111111"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2639
		when "101001001111" => B1 := "1111011"; B2 := "1111001"; B3 := "1011111"; B4 := "1101101"; 
		--2640
		when "101001010000" => B1 := "1111110"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2641
		when "101001010001" => B1 := "0110000"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2642
		when "101001010010" => B1 := "1101101"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2643
		when "101001010011" => B1 := "1111001"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2644
		when "101001010100" => B1 := "0110011"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2645
		when "101001010101" => B1 := "1011011"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2646
		when "101001010110" => B1 := "1011111"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2647
		when "101001010111" => B1 := "1110000"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2648
		when "101001011000" => B1 := "1111111"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2649
		when "101001011001" => B1 := "1111011"; B2 := "0110011"; B3 := "1011111"; B4 := "1101101"; 
		--2650
		when "101001011010" => B1 := "1111110"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2651
		when "101001011011" => B1 := "0110000"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2652
		when "101001011100" => B1 := "1101101"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2653
		when "101001011101" => B1 := "1111001"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2654
		when "101001011110" => B1 := "0110011"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2655
		when "101001011111" => B1 := "1011011"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2656
		when "101001100000" => B1 := "1011111"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2657
		when "101001100001" => B1 := "1110000"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2658
		when "101001100010" => B1 := "1111111"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2659
		when "101001100011" => B1 := "1111011"; B2 := "1011011"; B3 := "1011111"; B4 := "1101101"; 
		--2660
		when "101001100100" => B1 := "1111110"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2661
		when "101001100101" => B1 := "0110000"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2662
		when "101001100110" => B1 := "1101101"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2663
		when "101001100111" => B1 := "1111001"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2664
		when "101001101000" => B1 := "0110011"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2665
		when "101001101001" => B1 := "1011011"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2666
		when "101001101010" => B1 := "1011111"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2667
		when "101001101011" => B1 := "1110000"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2668
		when "101001101100" => B1 := "1111111"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2669
		when "101001101101" => B1 := "1111011"; B2 := "1011111"; B3 := "1011111"; B4 := "1101101"; 
		--2670
		when "101001101110" => B1 := "1111110"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2671
		when "101001101111" => B1 := "0110000"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2672
		when "101001110000" => B1 := "1101101"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2673
		when "101001110001" => B1 := "1111001"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2674
		when "101001110010" => B1 := "0110011"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2675
		when "101001110011" => B1 := "1011011"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2676
		when "101001110100" => B1 := "1011111"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2677
		when "101001110101" => B1 := "1110000"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2678
		when "101001110110" => B1 := "1111111"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2679
		when "101001110111" => B1 := "1111011"; B2 := "1110000"; B3 := "1011111"; B4 := "1101101"; 
		--2680
		when "101001111000" => B1 := "1111110"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2681
		when "101001111001" => B1 := "0110000"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2682
		when "101001111010" => B1 := "1101101"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2683
		when "101001111011" => B1 := "1111001"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2684
		when "101001111100" => B1 := "0110011"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2685
		when "101001111101" => B1 := "1011011"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2686
		when "101001111110" => B1 := "1011111"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2687
		when "101001111111" => B1 := "1110000"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2688
		when "101010000000" => B1 := "1111111"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2689
		when "101010000001" => B1 := "1111011"; B2 := "1111111"; B3 := "1011111"; B4 := "1101101"; 
		--2690
		when "101010000010" => B1 := "1111110"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2691
		when "101010000011" => B1 := "0110000"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2692
		when "101010000100" => B1 := "1101101"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2693
		when "101010000101" => B1 := "1111001"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2694
		when "101010000110" => B1 := "0110011"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2695
		when "101010000111" => B1 := "1011011"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2696
		when "101010001000" => B1 := "1011111"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2697
		when "101010001001" => B1 := "1110000"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2698
		when "101010001010" => B1 := "1111111"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2699
		when "101010001011" => B1 := "1111011"; B2 := "1111011"; B3 := "1011111"; B4 := "1101101"; 
		--2700
		when "101010001100" => B1 := "1111110"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2701
		when "101010001101" => B1 := "0110000"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2702
		when "101010001110" => B1 := "1101101"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2703
		when "101010001111" => B1 := "1111001"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2704
		when "101010010000" => B1 := "0110011"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2705
		when "101010010001" => B1 := "1011011"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2706
		when "101010010010" => B1 := "1011111"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2707
		when "101010010011" => B1 := "1110000"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2708
		when "101010010100" => B1 := "1111111"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2709
		when "101010010101" => B1 := "1111011"; B2 := "1111110"; B3 := "1110000"; B4 := "1101101"; 
		--2710
		when "101010010110" => B1 := "1111110"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2711
		when "101010010111" => B1 := "0110000"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2712
		when "101010011000" => B1 := "1101101"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2713
		when "101010011001" => B1 := "1111001"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2714
		when "101010011010" => B1 := "0110011"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2715
		when "101010011011" => B1 := "1011011"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2716
		when "101010011100" => B1 := "1011111"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2717
		when "101010011101" => B1 := "1110000"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2718
		when "101010011110" => B1 := "1111111"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2719
		when "101010011111" => B1 := "1111011"; B2 := "0110000"; B3 := "1110000"; B4 := "1101101"; 
		--2720
		when "101010100000" => B1 := "1111110"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2721
		when "101010100001" => B1 := "0110000"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2722
		when "101010100010" => B1 := "1101101"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2723
		when "101010100011" => B1 := "1111001"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2724
		when "101010100100" => B1 := "0110011"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2725
		when "101010100101" => B1 := "1011011"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2726
		when "101010100110" => B1 := "1011111"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2727
		when "101010100111" => B1 := "1110000"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2728
		when "101010101000" => B1 := "1111111"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2729
		when "101010101001" => B1 := "1111011"; B2 := "1101101"; B3 := "1110000"; B4 := "1101101"; 
		--2730
		when "101010101010" => B1 := "1111110"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2731
		when "101010101011" => B1 := "0110000"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2732
		when "101010101100" => B1 := "1101101"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2733
		when "101010101101" => B1 := "1111001"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2734
		when "101010101110" => B1 := "0110011"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2735
		when "101010101111" => B1 := "1011011"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2736
		when "101010110000" => B1 := "1011111"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2737
		when "101010110001" => B1 := "1110000"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2738
		when "101010110010" => B1 := "1111111"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2739
		when "101010110011" => B1 := "1111011"; B2 := "1111001"; B3 := "1110000"; B4 := "1101101"; 
		--2740
		when "101010110100" => B1 := "1111110"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2741
		when "101010110101" => B1 := "0110000"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2742
		when "101010110110" => B1 := "1101101"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2743
		when "101010110111" => B1 := "1111001"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2744
		when "101010111000" => B1 := "0110011"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2745
		when "101010111001" => B1 := "1011011"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2746
		when "101010111010" => B1 := "1011111"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2747
		when "101010111011" => B1 := "1110000"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2748
		when "101010111100" => B1 := "1111111"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2749
		when "101010111101" => B1 := "1111011"; B2 := "0110011"; B3 := "1110000"; B4 := "1101101"; 
		--2750
		when "101010111110" => B1 := "1111110"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2751
		when "101010111111" => B1 := "0110000"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2752
		when "101011000000" => B1 := "1101101"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2753
		when "101011000001" => B1 := "1111001"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2754
		when "101011000010" => B1 := "0110011"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2755
		when "101011000011" => B1 := "1011011"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2756
		when "101011000100" => B1 := "1011111"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2757
		when "101011000101" => B1 := "1110000"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2758
		when "101011000110" => B1 := "1111111"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2759
		when "101011000111" => B1 := "1111011"; B2 := "1011011"; B3 := "1110000"; B4 := "1101101"; 
		--2760
		when "101011001000" => B1 := "1111110"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2761
		when "101011001001" => B1 := "0110000"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2762
		when "101011001010" => B1 := "1101101"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2763
		when "101011001011" => B1 := "1111001"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2764
		when "101011001100" => B1 := "0110011"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2765
		when "101011001101" => B1 := "1011011"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2766
		when "101011001110" => B1 := "1011111"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2767
		when "101011001111" => B1 := "1110000"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2768
		when "101011010000" => B1 := "1111111"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2769
		when "101011010001" => B1 := "1111011"; B2 := "1011111"; B3 := "1110000"; B4 := "1101101"; 
		--2770
		when "101011010010" => B1 := "1111110"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2771
		when "101011010011" => B1 := "0110000"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2772
		when "101011010100" => B1 := "1101101"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2773
		when "101011010101" => B1 := "1111001"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2774
		when "101011010110" => B1 := "0110011"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2775
		when "101011010111" => B1 := "1011011"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2776
		when "101011011000" => B1 := "1011111"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2777
		when "101011011001" => B1 := "1110000"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2778
		when "101011011010" => B1 := "1111111"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2779
		when "101011011011" => B1 := "1111011"; B2 := "1110000"; B3 := "1110000"; B4 := "1101101"; 
		--2780
		when "101011011100" => B1 := "1111110"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2781
		when "101011011101" => B1 := "0110000"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2782
		when "101011011110" => B1 := "1101101"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2783
		when "101011011111" => B1 := "1111001"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2784
		when "101011100000" => B1 := "0110011"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2785
		when "101011100001" => B1 := "1011011"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2786
		when "101011100010" => B1 := "1011111"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2787
		when "101011100011" => B1 := "1110000"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2788
		when "101011100100" => B1 := "1111111"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2789
		when "101011100101" => B1 := "1111011"; B2 := "1111111"; B3 := "1110000"; B4 := "1101101"; 
		--2790
		when "101011100110" => B1 := "1111110"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2791
		when "101011100111" => B1 := "0110000"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2792
		when "101011101000" => B1 := "1101101"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2793
		when "101011101001" => B1 := "1111001"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2794
		when "101011101010" => B1 := "0110011"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2795
		when "101011101011" => B1 := "1011011"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2796
		when "101011101100" => B1 := "1011111"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2797
		when "101011101101" => B1 := "1110000"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2798
		when "101011101110" => B1 := "1111111"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2799
		when "101011101111" => B1 := "1111011"; B2 := "1111011"; B3 := "1110000"; B4 := "1101101"; 
		--2800
		when "101011110000" => B1 := "1111110"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2801
		when "101011110001" => B1 := "0110000"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2802
		when "101011110010" => B1 := "1101101"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2803
		when "101011110011" => B1 := "1111001"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2804
		when "101011110100" => B1 := "0110011"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2805
		when "101011110101" => B1 := "1011011"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2806
		when "101011110110" => B1 := "1011111"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2807
		when "101011110111" => B1 := "1110000"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2808
		when "101011111000" => B1 := "1111111"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2809
		when "101011111001" => B1 := "1111011"; B2 := "1111110"; B3 := "1111111"; B4 := "1101101"; 
		--2810
		when "101011111010" => B1 := "1111110"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2811
		when "101011111011" => B1 := "0110000"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2812
		when "101011111100" => B1 := "1101101"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2813
		when "101011111101" => B1 := "1111001"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2814
		when "101011111110" => B1 := "0110011"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2815
		when "101011111111" => B1 := "1011011"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2816
		when "101100000000" => B1 := "1011111"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2817
		when "101100000001" => B1 := "1110000"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2818
		when "101100000010" => B1 := "1111111"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2819
		when "101100000011" => B1 := "1111011"; B2 := "0110000"; B3 := "1111111"; B4 := "1101101"; 
		--2820
		when "101100000100" => B1 := "1111110"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2821
		when "101100000101" => B1 := "0110000"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2822
		when "101100000110" => B1 := "1101101"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2823
		when "101100000111" => B1 := "1111001"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2824
		when "101100001000" => B1 := "0110011"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2825
		when "101100001001" => B1 := "1011011"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2826
		when "101100001010" => B1 := "1011111"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2827
		when "101100001011" => B1 := "1110000"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2828
		when "101100001100" => B1 := "1111111"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2829
		when "101100001101" => B1 := "1111011"; B2 := "1101101"; B3 := "1111111"; B4 := "1101101"; 
		--2830
		when "101100001110" => B1 := "1111110"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2831
		when "101100001111" => B1 := "0110000"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2832
		when "101100010000" => B1 := "1101101"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2833
		when "101100010001" => B1 := "1111001"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2834
		when "101100010010" => B1 := "0110011"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2835
		when "101100010011" => B1 := "1011011"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2836
		when "101100010100" => B1 := "1011111"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2837
		when "101100010101" => B1 := "1110000"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2838
		when "101100010110" => B1 := "1111111"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2839
		when "101100010111" => B1 := "1111011"; B2 := "1111001"; B3 := "1111111"; B4 := "1101101"; 
		--2840
		when "101100011000" => B1 := "1111110"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2841
		when "101100011001" => B1 := "0110000"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2842
		when "101100011010" => B1 := "1101101"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2843
		when "101100011011" => B1 := "1111001"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2844
		when "101100011100" => B1 := "0110011"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2845
		when "101100011101" => B1 := "1011011"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2846
		when "101100011110" => B1 := "1011111"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2847
		when "101100011111" => B1 := "1110000"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2848
		when "101100100000" => B1 := "1111111"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2849
		when "101100100001" => B1 := "1111011"; B2 := "0110011"; B3 := "1111111"; B4 := "1101101"; 
		--2850
		when "101100100010" => B1 := "1111110"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2851
		when "101100100011" => B1 := "0110000"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2852
		when "101100100100" => B1 := "1101101"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2853
		when "101100100101" => B1 := "1111001"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2854
		when "101100100110" => B1 := "0110011"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2855
		when "101100100111" => B1 := "1011011"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2856
		when "101100101000" => B1 := "1011111"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2857
		when "101100101001" => B1 := "1110000"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2858
		when "101100101010" => B1 := "1111111"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2859
		when "101100101011" => B1 := "1111011"; B2 := "1011011"; B3 := "1111111"; B4 := "1101101"; 
		--2860
		when "101100101100" => B1 := "1111110"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2861
		when "101100101101" => B1 := "0110000"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2862
		when "101100101110" => B1 := "1101101"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2863
		when "101100101111" => B1 := "1111001"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2864
		when "101100110000" => B1 := "0110011"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2865
		when "101100110001" => B1 := "1011011"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2866
		when "101100110010" => B1 := "1011111"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2867
		when "101100110011" => B1 := "1110000"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2868
		when "101100110100" => B1 := "1111111"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2869
		when "101100110101" => B1 := "1111011"; B2 := "1011111"; B3 := "1111111"; B4 := "1101101"; 
		--2870
		when "101100110110" => B1 := "1111110"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2871
		when "101100110111" => B1 := "0110000"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2872
		when "101100111000" => B1 := "1101101"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2873
		when "101100111001" => B1 := "1111001"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2874
		when "101100111010" => B1 := "0110011"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2875
		when "101100111011" => B1 := "1011011"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2876
		when "101100111100" => B1 := "1011111"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2877
		when "101100111101" => B1 := "1110000"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2878
		when "101100111110" => B1 := "1111111"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2879
		when "101100111111" => B1 := "1111011"; B2 := "1110000"; B3 := "1111111"; B4 := "1101101"; 
		--2880
		when "101101000000" => B1 := "1111110"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2881
		when "101101000001" => B1 := "0110000"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2882
		when "101101000010" => B1 := "1101101"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2883
		when "101101000011" => B1 := "1111001"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2884
		when "101101000100" => B1 := "0110011"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2885
		when "101101000101" => B1 := "1011011"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2886
		when "101101000110" => B1 := "1011111"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2887
		when "101101000111" => B1 := "1110000"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2888
		when "101101001000" => B1 := "1111111"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2889
		when "101101001001" => B1 := "1111011"; B2 := "1111111"; B3 := "1111111"; B4 := "1101101"; 
		--2890
		when "101101001010" => B1 := "1111110"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2891
		when "101101001011" => B1 := "0110000"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2892
		when "101101001100" => B1 := "1101101"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2893
		when "101101001101" => B1 := "1111001"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2894
		when "101101001110" => B1 := "0110011"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2895
		when "101101001111" => B1 := "1011011"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2896
		when "101101010000" => B1 := "1011111"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2897
		when "101101010001" => B1 := "1110000"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2898
		when "101101010010" => B1 := "1111111"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2899
		when "101101010011" => B1 := "1111011"; B2 := "1111011"; B3 := "1111111"; B4 := "1101101"; 
		--2900
		when "101101010100" => B1 := "1111110"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2901
		when "101101010101" => B1 := "0110000"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2902
		when "101101010110" => B1 := "1101101"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2903
		when "101101010111" => B1 := "1111001"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2904
		when "101101011000" => B1 := "0110011"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2905
		when "101101011001" => B1 := "1011011"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2906
		when "101101011010" => B1 := "1011111"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2907
		when "101101011011" => B1 := "1110000"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2908
		when "101101011100" => B1 := "1111111"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2909
		when "101101011101" => B1 := "1111011"; B2 := "1111110"; B3 := "1111011"; B4 := "1101101"; 
		--2910
		when "101101011110" => B1 := "1111110"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2911
		when "101101011111" => B1 := "0110000"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2912
		when "101101100000" => B1 := "1101101"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2913
		when "101101100001" => B1 := "1111001"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2914
		when "101101100010" => B1 := "0110011"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2915
		when "101101100011" => B1 := "1011011"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2916
		when "101101100100" => B1 := "1011111"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2917
		when "101101100101" => B1 := "1110000"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2918
		when "101101100110" => B1 := "1111111"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2919
		when "101101100111" => B1 := "1111011"; B2 := "0110000"; B3 := "1111011"; B4 := "1101101"; 
		--2920
		when "101101101000" => B1 := "1111110"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2921
		when "101101101001" => B1 := "0110000"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2922
		when "101101101010" => B1 := "1101101"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2923
		when "101101101011" => B1 := "1111001"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2924
		when "101101101100" => B1 := "0110011"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2925
		when "101101101101" => B1 := "1011011"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2926
		when "101101101110" => B1 := "1011111"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2927
		when "101101101111" => B1 := "1110000"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2928
		when "101101110000" => B1 := "1111111"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2929
		when "101101110001" => B1 := "1111011"; B2 := "1101101"; B3 := "1111011"; B4 := "1101101"; 
		--2930
		when "101101110010" => B1 := "1111110"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2931
		when "101101110011" => B1 := "0110000"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2932
		when "101101110100" => B1 := "1101101"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2933
		when "101101110101" => B1 := "1111001"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2934
		when "101101110110" => B1 := "0110011"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2935
		when "101101110111" => B1 := "1011011"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2936
		when "101101111000" => B1 := "1011111"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2937
		when "101101111001" => B1 := "1110000"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2938
		when "101101111010" => B1 := "1111111"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2939
		when "101101111011" => B1 := "1111011"; B2 := "1111001"; B3 := "1111011"; B4 := "1101101"; 
		--2940
		when "101101111100" => B1 := "1111110"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2941
		when "101101111101" => B1 := "0110000"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2942
		when "101101111110" => B1 := "1101101"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2943
		when "101101111111" => B1 := "1111001"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2944
		when "101110000000" => B1 := "0110011"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2945
		when "101110000001" => B1 := "1011011"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2946
		when "101110000010" => B1 := "1011111"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2947
		when "101110000011" => B1 := "1110000"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2948
		when "101110000100" => B1 := "1111111"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2949
		when "101110000101" => B1 := "1111011"; B2 := "0110011"; B3 := "1111011"; B4 := "1101101"; 
		--2950
		when "101110000110" => B1 := "1111110"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2951
		when "101110000111" => B1 := "0110000"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2952
		when "101110001000" => B1 := "1101101"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2953
		when "101110001001" => B1 := "1111001"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2954
		when "101110001010" => B1 := "0110011"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2955
		when "101110001011" => B1 := "1011011"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2956
		when "101110001100" => B1 := "1011111"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2957
		when "101110001101" => B1 := "1110000"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2958
		when "101110001110" => B1 := "1111111"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2959
		when "101110001111" => B1 := "1111011"; B2 := "1011011"; B3 := "1111011"; B4 := "1101101"; 
		--2960
		when "101110010000" => B1 := "1111110"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2961
		when "101110010001" => B1 := "0110000"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2962
		when "101110010010" => B1 := "1101101"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2963
		when "101110010011" => B1 := "1111001"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2964
		when "101110010100" => B1 := "0110011"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2965
		when "101110010101" => B1 := "1011011"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2966
		when "101110010110" => B1 := "1011111"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2967
		when "101110010111" => B1 := "1110000"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2968
		when "101110011000" => B1 := "1111111"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2969
		when "101110011001" => B1 := "1111011"; B2 := "1011111"; B3 := "1111011"; B4 := "1101101"; 
		--2970
		when "101110011010" => B1 := "1111110"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2971
		when "101110011011" => B1 := "0110000"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2972
		when "101110011100" => B1 := "1101101"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2973
		when "101110011101" => B1 := "1111001"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2974
		when "101110011110" => B1 := "0110011"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2975
		when "101110011111" => B1 := "1011011"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2976
		when "101110100000" => B1 := "1011111"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2977
		when "101110100001" => B1 := "1110000"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2978
		when "101110100010" => B1 := "1111111"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2979
		when "101110100011" => B1 := "1111011"; B2 := "1110000"; B3 := "1111011"; B4 := "1101101"; 
		--2980
		when "101110100100" => B1 := "1111110"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2981
		when "101110100101" => B1 := "0110000"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2982
		when "101110100110" => B1 := "1101101"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2983
		when "101110100111" => B1 := "1111001"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2984
		when "101110101000" => B1 := "0110011"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2985
		when "101110101001" => B1 := "1011011"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2986
		when "101110101010" => B1 := "1011111"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2987
		when "101110101011" => B1 := "1110000"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2988
		when "101110101100" => B1 := "1111111"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2989
		when "101110101101" => B1 := "1111011"; B2 := "1111111"; B3 := "1111011"; B4 := "1101101"; 
		--2990
		when "101110101110" => B1 := "1111110"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--2991
		when "101110101111" => B1 := "0110000"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--2992
		when "101110110000" => B1 := "1101101"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--2993
		when "101110110001" => B1 := "1111001"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--2994
		when "101110110010" => B1 := "0110011"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--2995
		when "101110110011" => B1 := "1011011"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--2996
		when "101110110100" => B1 := "1011111"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--2997
		when "101110110101" => B1 := "1110000"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--2998
		when "101110110110" => B1 := "1111111"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--2999
		when "101110110111" => B1 := "1111011"; B2 := "1111011"; B3 := "1111011"; B4 := "1101101"; 
		--3000
		when "101110111000" => B1 := "1111110"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3001
		when "101110111001" => B1 := "0110000"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3002
		when "101110111010" => B1 := "1101101"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3003
		when "101110111011" => B1 := "1111001"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3004
		when "101110111100" => B1 := "0110011"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3005
		when "101110111101" => B1 := "1011011"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3006
		when "101110111110" => B1 := "1011111"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3007
		when "101110111111" => B1 := "1110000"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3008
		when "101111000000" => B1 := "1111111"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3009
		when "101111000001" => B1 := "1111011"; B2 := "1111110"; B3 := "1111110"; B4 := "1111001"; 
		--3010
		when "101111000010" => B1 := "1111110"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3011
		when "101111000011" => B1 := "0110000"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3012
		when "101111000100" => B1 := "1101101"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3013
		when "101111000101" => B1 := "1111001"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3014
		when "101111000110" => B1 := "0110011"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3015
		when "101111000111" => B1 := "1011011"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3016
		when "101111001000" => B1 := "1011111"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3017
		when "101111001001" => B1 := "1110000"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3018
		when "101111001010" => B1 := "1111111"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3019
		when "101111001011" => B1 := "1111011"; B2 := "0110000"; B3 := "1111110"; B4 := "1111001"; 
		--3020
		when "101111001100" => B1 := "1111110"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3021
		when "101111001101" => B1 := "0110000"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3022
		when "101111001110" => B1 := "1101101"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3023
		when "101111001111" => B1 := "1111001"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3024
		when "101111010000" => B1 := "0110011"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3025
		when "101111010001" => B1 := "1011011"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3026
		when "101111010010" => B1 := "1011111"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3027
		when "101111010011" => B1 := "1110000"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3028
		when "101111010100" => B1 := "1111111"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3029
		when "101111010101" => B1 := "1111011"; B2 := "1101101"; B3 := "1111110"; B4 := "1111001"; 
		--3030
		when "101111010110" => B1 := "1111110"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3031
		when "101111010111" => B1 := "0110000"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3032
		when "101111011000" => B1 := "1101101"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3033
		when "101111011001" => B1 := "1111001"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3034
		when "101111011010" => B1 := "0110011"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3035
		when "101111011011" => B1 := "1011011"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3036
		when "101111011100" => B1 := "1011111"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3037
		when "101111011101" => B1 := "1110000"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3038
		when "101111011110" => B1 := "1111111"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3039
		when "101111011111" => B1 := "1111011"; B2 := "1111001"; B3 := "1111110"; B4 := "1111001"; 
		--3040
		when "101111100000" => B1 := "1111110"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3041
		when "101111100001" => B1 := "0110000"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3042
		when "101111100010" => B1 := "1101101"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3043
		when "101111100011" => B1 := "1111001"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3044
		when "101111100100" => B1 := "0110011"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3045
		when "101111100101" => B1 := "1011011"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3046
		when "101111100110" => B1 := "1011111"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3047
		when "101111100111" => B1 := "1110000"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3048
		when "101111101000" => B1 := "1111111"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3049
		when "101111101001" => B1 := "1111011"; B2 := "0110011"; B3 := "1111110"; B4 := "1111001"; 
		--3050
		when "101111101010" => B1 := "1111110"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3051
		when "101111101011" => B1 := "0110000"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3052
		when "101111101100" => B1 := "1101101"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3053
		when "101111101101" => B1 := "1111001"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3054
		when "101111101110" => B1 := "0110011"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3055
		when "101111101111" => B1 := "1011011"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3056
		when "101111110000" => B1 := "1011111"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3057
		when "101111110001" => B1 := "1110000"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3058
		when "101111110010" => B1 := "1111111"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3059
		when "101111110011" => B1 := "1111011"; B2 := "1011011"; B3 := "1111110"; B4 := "1111001"; 
		--3060
		when "101111110100" => B1 := "1111110"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3061
		when "101111110101" => B1 := "0110000"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3062
		when "101111110110" => B1 := "1101101"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3063
		when "101111110111" => B1 := "1111001"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3064
		when "101111111000" => B1 := "0110011"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3065
		when "101111111001" => B1 := "1011011"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3066
		when "101111111010" => B1 := "1011111"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3067
		when "101111111011" => B1 := "1110000"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3068
		when "101111111100" => B1 := "1111111"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3069
		when "101111111101" => B1 := "1111011"; B2 := "1011111"; B3 := "1111110"; B4 := "1111001"; 
		--3070
		when "101111111110" => B1 := "1111110"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3071
		when "101111111111" => B1 := "0110000"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3072
		when "110000000000" => B1 := "1101101"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3073
		when "110000000001" => B1 := "1111001"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3074
		when "110000000010" => B1 := "0110011"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3075
		when "110000000011" => B1 := "1011011"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3076
		when "110000000100" => B1 := "1011111"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3077
		when "110000000101" => B1 := "1110000"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3078
		when "110000000110" => B1 := "1111111"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3079
		when "110000000111" => B1 := "1111011"; B2 := "1110000"; B3 := "1111110"; B4 := "1111001"; 
		--3080
		when "110000001000" => B1 := "1111110"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3081
		when "110000001001" => B1 := "0110000"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3082
		when "110000001010" => B1 := "1101101"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3083
		when "110000001011" => B1 := "1111001"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3084
		when "110000001100" => B1 := "0110011"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3085
		when "110000001101" => B1 := "1011011"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3086
		when "110000001110" => B1 := "1011111"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3087
		when "110000001111" => B1 := "1110000"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3088
		when "110000010000" => B1 := "1111111"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3089
		when "110000010001" => B1 := "1111011"; B2 := "1111111"; B3 := "1111110"; B4 := "1111001"; 
		--3090
		when "110000010010" => B1 := "1111110"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3091
		when "110000010011" => B1 := "0110000"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3092
		when "110000010100" => B1 := "1101101"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3093
		when "110000010101" => B1 := "1111001"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3094
		when "110000010110" => B1 := "0110011"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3095
		when "110000010111" => B1 := "1011011"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3096
		when "110000011000" => B1 := "1011111"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3097
		when "110000011001" => B1 := "1110000"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3098
		when "110000011010" => B1 := "1111111"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3099
		when "110000011011" => B1 := "1111011"; B2 := "1111011"; B3 := "1111110"; B4 := "1111001"; 
		--3100
		when "110000011100" => B1 := "1111110"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3101
		when "110000011101" => B1 := "0110000"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3102
		when "110000011110" => B1 := "1101101"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3103
		when "110000011111" => B1 := "1111001"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3104
		when "110000100000" => B1 := "0110011"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3105
		when "110000100001" => B1 := "1011011"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3106
		when "110000100010" => B1 := "1011111"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3107
		when "110000100011" => B1 := "1110000"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3108
		when "110000100100" => B1 := "1111111"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3109
		when "110000100101" => B1 := "1111011"; B2 := "1111110"; B3 := "0110000"; B4 := "1111001"; 
		--3110
		when "110000100110" => B1 := "1111110"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3111
		when "110000100111" => B1 := "0110000"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3112
		when "110000101000" => B1 := "1101101"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3113
		when "110000101001" => B1 := "1111001"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3114
		when "110000101010" => B1 := "0110011"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3115
		when "110000101011" => B1 := "1011011"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3116
		when "110000101100" => B1 := "1011111"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3117
		when "110000101101" => B1 := "1110000"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3118
		when "110000101110" => B1 := "1111111"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3119
		when "110000101111" => B1 := "1111011"; B2 := "0110000"; B3 := "0110000"; B4 := "1111001"; 
		--3120
		when "110000110000" => B1 := "1111110"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3121
		when "110000110001" => B1 := "0110000"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3122
		when "110000110010" => B1 := "1101101"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3123
		when "110000110011" => B1 := "1111001"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3124
		when "110000110100" => B1 := "0110011"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3125
		when "110000110101" => B1 := "1011011"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3126
		when "110000110110" => B1 := "1011111"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3127
		when "110000110111" => B1 := "1110000"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3128
		when "110000111000" => B1 := "1111111"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3129
		when "110000111001" => B1 := "1111011"; B2 := "1101101"; B3 := "0110000"; B4 := "1111001"; 
		--3130
		when "110000111010" => B1 := "1111110"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3131
		when "110000111011" => B1 := "0110000"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3132
		when "110000111100" => B1 := "1101101"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3133
		when "110000111101" => B1 := "1111001"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3134
		when "110000111110" => B1 := "0110011"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3135
		when "110000111111" => B1 := "1011011"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3136
		when "110001000000" => B1 := "1011111"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3137
		when "110001000001" => B1 := "1110000"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3138
		when "110001000010" => B1 := "1111111"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3139
		when "110001000011" => B1 := "1111011"; B2 := "1111001"; B3 := "0110000"; B4 := "1111001"; 
		--3140
		when "110001000100" => B1 := "1111110"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3141
		when "110001000101" => B1 := "0110000"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3142
		when "110001000110" => B1 := "1101101"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3143
		when "110001000111" => B1 := "1111001"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3144
		when "110001001000" => B1 := "0110011"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3145
		when "110001001001" => B1 := "1011011"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3146
		when "110001001010" => B1 := "1011111"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3147
		when "110001001011" => B1 := "1110000"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3148
		when "110001001100" => B1 := "1111111"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3149
		when "110001001101" => B1 := "1111011"; B2 := "0110011"; B3 := "0110000"; B4 := "1111001"; 
		--3150
		when "110001001110" => B1 := "1111110"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3151
		when "110001001111" => B1 := "0110000"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3152
		when "110001010000" => B1 := "1101101"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3153
		when "110001010001" => B1 := "1111001"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3154
		when "110001010010" => B1 := "0110011"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3155
		when "110001010011" => B1 := "1011011"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3156
		when "110001010100" => B1 := "1011111"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3157
		when "110001010101" => B1 := "1110000"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3158
		when "110001010110" => B1 := "1111111"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3159
		when "110001010111" => B1 := "1111011"; B2 := "1011011"; B3 := "0110000"; B4 := "1111001"; 
		--3160
		when "110001011000" => B1 := "1111110"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3161
		when "110001011001" => B1 := "0110000"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3162
		when "110001011010" => B1 := "1101101"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3163
		when "110001011011" => B1 := "1111001"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3164
		when "110001011100" => B1 := "0110011"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3165
		when "110001011101" => B1 := "1011011"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3166
		when "110001011110" => B1 := "1011111"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3167
		when "110001011111" => B1 := "1110000"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3168
		when "110001100000" => B1 := "1111111"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3169
		when "110001100001" => B1 := "1111011"; B2 := "1011111"; B3 := "0110000"; B4 := "1111001"; 
		--3170
		when "110001100010" => B1 := "1111110"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3171
		when "110001100011" => B1 := "0110000"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3172
		when "110001100100" => B1 := "1101101"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3173
		when "110001100101" => B1 := "1111001"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3174
		when "110001100110" => B1 := "0110011"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3175
		when "110001100111" => B1 := "1011011"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3176
		when "110001101000" => B1 := "1011111"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3177
		when "110001101001" => B1 := "1110000"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3178
		when "110001101010" => B1 := "1111111"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3179
		when "110001101011" => B1 := "1111011"; B2 := "1110000"; B3 := "0110000"; B4 := "1111001"; 
		--3180
		when "110001101100" => B1 := "1111110"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3181
		when "110001101101" => B1 := "0110000"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3182
		when "110001101110" => B1 := "1101101"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3183
		when "110001101111" => B1 := "1111001"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3184
		when "110001110000" => B1 := "0110011"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3185
		when "110001110001" => B1 := "1011011"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3186
		when "110001110010" => B1 := "1011111"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3187
		when "110001110011" => B1 := "1110000"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3188
		when "110001110100" => B1 := "1111111"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3189
		when "110001110101" => B1 := "1111011"; B2 := "1111111"; B3 := "0110000"; B4 := "1111001"; 
		--3190
		when "110001110110" => B1 := "1111110"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3191
		when "110001110111" => B1 := "0110000"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3192
		when "110001111000" => B1 := "1101101"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3193
		when "110001111001" => B1 := "1111001"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3194
		when "110001111010" => B1 := "0110011"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3195
		when "110001111011" => B1 := "1011011"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3196
		when "110001111100" => B1 := "1011111"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3197
		when "110001111101" => B1 := "1110000"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3198
		when "110001111110" => B1 := "1111111"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3199
		when "110001111111" => B1 := "1111011"; B2 := "1111011"; B3 := "0110000"; B4 := "1111001"; 
		--3200
		when "110010000000" => B1 := "1111110"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3201
		when "110010000001" => B1 := "0110000"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3202
		when "110010000010" => B1 := "1101101"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3203
		when "110010000011" => B1 := "1111001"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3204
		when "110010000100" => B1 := "0110011"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3205
		when "110010000101" => B1 := "1011011"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3206
		when "110010000110" => B1 := "1011111"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3207
		when "110010000111" => B1 := "1110000"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3208
		when "110010001000" => B1 := "1111111"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3209
		when "110010001001" => B1 := "1111011"; B2 := "1111110"; B3 := "1101101"; B4 := "1111001"; 
		--3210
		when "110010001010" => B1 := "1111110"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3211
		when "110010001011" => B1 := "0110000"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3212
		when "110010001100" => B1 := "1101101"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3213
		when "110010001101" => B1 := "1111001"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3214
		when "110010001110" => B1 := "0110011"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3215
		when "110010001111" => B1 := "1011011"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3216
		when "110010010000" => B1 := "1011111"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3217
		when "110010010001" => B1 := "1110000"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3218
		when "110010010010" => B1 := "1111111"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3219
		when "110010010011" => B1 := "1111011"; B2 := "0110000"; B3 := "1101101"; B4 := "1111001"; 
		--3220
		when "110010010100" => B1 := "1111110"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3221
		when "110010010101" => B1 := "0110000"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3222
		when "110010010110" => B1 := "1101101"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3223
		when "110010010111" => B1 := "1111001"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3224
		when "110010011000" => B1 := "0110011"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3225
		when "110010011001" => B1 := "1011011"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3226
		when "110010011010" => B1 := "1011111"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3227
		when "110010011011" => B1 := "1110000"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3228
		when "110010011100" => B1 := "1111111"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3229
		when "110010011101" => B1 := "1111011"; B2 := "1101101"; B3 := "1101101"; B4 := "1111001"; 
		--3230
		when "110010011110" => B1 := "1111110"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3231
		when "110010011111" => B1 := "0110000"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3232
		when "110010100000" => B1 := "1101101"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3233
		when "110010100001" => B1 := "1111001"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3234
		when "110010100010" => B1 := "0110011"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3235
		when "110010100011" => B1 := "1011011"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3236
		when "110010100100" => B1 := "1011111"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3237
		when "110010100101" => B1 := "1110000"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3238
		when "110010100110" => B1 := "1111111"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3239
		when "110010100111" => B1 := "1111011"; B2 := "1111001"; B3 := "1101101"; B4 := "1111001"; 
		--3240
		when "110010101000" => B1 := "1111110"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3241
		when "110010101001" => B1 := "0110000"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3242
		when "110010101010" => B1 := "1101101"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3243
		when "110010101011" => B1 := "1111001"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3244
		when "110010101100" => B1 := "0110011"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3245
		when "110010101101" => B1 := "1011011"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3246
		when "110010101110" => B1 := "1011111"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3247
		when "110010101111" => B1 := "1110000"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3248
		when "110010110000" => B1 := "1111111"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3249
		when "110010110001" => B1 := "1111011"; B2 := "0110011"; B3 := "1101101"; B4 := "1111001"; 
		--3250
		when "110010110010" => B1 := "1111110"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3251
		when "110010110011" => B1 := "0110000"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3252
		when "110010110100" => B1 := "1101101"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3253
		when "110010110101" => B1 := "1111001"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3254
		when "110010110110" => B1 := "0110011"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3255
		when "110010110111" => B1 := "1011011"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3256
		when "110010111000" => B1 := "1011111"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3257
		when "110010111001" => B1 := "1110000"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3258
		when "110010111010" => B1 := "1111111"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3259
		when "110010111011" => B1 := "1111011"; B2 := "1011011"; B3 := "1101101"; B4 := "1111001"; 
		--3260
		when "110010111100" => B1 := "1111110"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3261
		when "110010111101" => B1 := "0110000"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3262
		when "110010111110" => B1 := "1101101"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3263
		when "110010111111" => B1 := "1111001"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3264
		when "110011000000" => B1 := "0110011"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3265
		when "110011000001" => B1 := "1011011"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3266
		when "110011000010" => B1 := "1011111"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3267
		when "110011000011" => B1 := "1110000"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3268
		when "110011000100" => B1 := "1111111"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3269
		when "110011000101" => B1 := "1111011"; B2 := "1011111"; B3 := "1101101"; B4 := "1111001"; 
		--3270
		when "110011000110" => B1 := "1111110"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3271
		when "110011000111" => B1 := "0110000"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3272
		when "110011001000" => B1 := "1101101"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3273
		when "110011001001" => B1 := "1111001"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3274
		when "110011001010" => B1 := "0110011"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3275
		when "110011001011" => B1 := "1011011"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3276
		when "110011001100" => B1 := "1011111"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3277
		when "110011001101" => B1 := "1110000"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3278
		when "110011001110" => B1 := "1111111"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3279
		when "110011001111" => B1 := "1111011"; B2 := "1110000"; B3 := "1101101"; B4 := "1111001"; 
		--3280
		when "110011010000" => B1 := "1111110"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3281
		when "110011010001" => B1 := "0110000"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3282
		when "110011010010" => B1 := "1101101"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3283
		when "110011010011" => B1 := "1111001"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3284
		when "110011010100" => B1 := "0110011"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3285
		when "110011010101" => B1 := "1011011"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3286
		when "110011010110" => B1 := "1011111"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3287
		when "110011010111" => B1 := "1110000"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3288
		when "110011011000" => B1 := "1111111"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3289
		when "110011011001" => B1 := "1111011"; B2 := "1111111"; B3 := "1101101"; B4 := "1111001"; 
		--3290
		when "110011011010" => B1 := "1111110"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3291
		when "110011011011" => B1 := "0110000"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3292
		when "110011011100" => B1 := "1101101"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3293
		when "110011011101" => B1 := "1111001"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3294
		when "110011011110" => B1 := "0110011"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3295
		when "110011011111" => B1 := "1011011"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3296
		when "110011100000" => B1 := "1011111"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3297
		when "110011100001" => B1 := "1110000"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3298
		when "110011100010" => B1 := "1111111"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3299
		when "110011100011" => B1 := "1111011"; B2 := "1111011"; B3 := "1101101"; B4 := "1111001"; 
		--3300
		when "110011100100" => B1 := "1111110"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3301
		when "110011100101" => B1 := "0110000"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3302
		when "110011100110" => B1 := "1101101"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3303
		when "110011100111" => B1 := "1111001"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3304
		when "110011101000" => B1 := "0110011"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3305
		when "110011101001" => B1 := "1011011"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3306
		when "110011101010" => B1 := "1011111"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3307
		when "110011101011" => B1 := "1110000"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3308
		when "110011101100" => B1 := "1111111"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3309
		when "110011101101" => B1 := "1111011"; B2 := "1111110"; B3 := "1111001"; B4 := "1111001"; 
		--3310
		when "110011101110" => B1 := "1111110"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3311
		when "110011101111" => B1 := "0110000"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3312
		when "110011110000" => B1 := "1101101"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3313
		when "110011110001" => B1 := "1111001"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3314
		when "110011110010" => B1 := "0110011"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3315
		when "110011110011" => B1 := "1011011"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3316
		when "110011110100" => B1 := "1011111"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3317
		when "110011110101" => B1 := "1110000"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3318
		when "110011110110" => B1 := "1111111"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3319
		when "110011110111" => B1 := "1111011"; B2 := "0110000"; B3 := "1111001"; B4 := "1111001"; 
		--3320
		when "110011111000" => B1 := "1111110"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3321
		when "110011111001" => B1 := "0110000"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3322
		when "110011111010" => B1 := "1101101"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3323
		when "110011111011" => B1 := "1111001"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3324
		when "110011111100" => B1 := "0110011"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3325
		when "110011111101" => B1 := "1011011"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3326
		when "110011111110" => B1 := "1011111"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3327
		when "110011111111" => B1 := "1110000"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3328
		when "110100000000" => B1 := "1111111"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3329
		when "110100000001" => B1 := "1111011"; B2 := "1101101"; B3 := "1111001"; B4 := "1111001"; 
		--3330
		when "110100000010" => B1 := "1111110"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3331
		when "110100000011" => B1 := "0110000"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3332
		when "110100000100" => B1 := "1101101"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3333
		when "110100000101" => B1 := "1111001"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3334
		when "110100000110" => B1 := "0110011"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3335
		when "110100000111" => B1 := "1011011"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3336
		when "110100001000" => B1 := "1011111"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3337
		when "110100001001" => B1 := "1110000"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3338
		when "110100001010" => B1 := "1111111"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3339
		when "110100001011" => B1 := "1111011"; B2 := "1111001"; B3 := "1111001"; B4 := "1111001"; 
		--3340
		when "110100001100" => B1 := "1111110"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3341
		when "110100001101" => B1 := "0110000"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3342
		when "110100001110" => B1 := "1101101"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3343
		when "110100001111" => B1 := "1111001"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3344
		when "110100010000" => B1 := "0110011"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3345
		when "110100010001" => B1 := "1011011"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3346
		when "110100010010" => B1 := "1011111"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3347
		when "110100010011" => B1 := "1110000"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3348
		when "110100010100" => B1 := "1111111"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3349
		when "110100010101" => B1 := "1111011"; B2 := "0110011"; B3 := "1111001"; B4 := "1111001"; 
		--3350
		when "110100010110" => B1 := "1111110"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3351
		when "110100010111" => B1 := "0110000"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3352
		when "110100011000" => B1 := "1101101"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3353
		when "110100011001" => B1 := "1111001"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3354
		when "110100011010" => B1 := "0110011"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3355
		when "110100011011" => B1 := "1011011"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3356
		when "110100011100" => B1 := "1011111"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3357
		when "110100011101" => B1 := "1110000"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3358
		when "110100011110" => B1 := "1111111"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3359
		when "110100011111" => B1 := "1111011"; B2 := "1011011"; B3 := "1111001"; B4 := "1111001"; 
		--3360
		when "110100100000" => B1 := "1111110"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3361
		when "110100100001" => B1 := "0110000"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3362
		when "110100100010" => B1 := "1101101"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3363
		when "110100100011" => B1 := "1111001"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3364
		when "110100100100" => B1 := "0110011"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3365
		when "110100100101" => B1 := "1011011"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3366
		when "110100100110" => B1 := "1011111"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3367
		when "110100100111" => B1 := "1110000"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3368
		when "110100101000" => B1 := "1111111"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3369
		when "110100101001" => B1 := "1111011"; B2 := "1011111"; B3 := "1111001"; B4 := "1111001"; 
		--3370
		when "110100101010" => B1 := "1111110"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3371
		when "110100101011" => B1 := "0110000"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3372
		when "110100101100" => B1 := "1101101"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3373
		when "110100101101" => B1 := "1111001"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3374
		when "110100101110" => B1 := "0110011"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3375
		when "110100101111" => B1 := "1011011"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3376
		when "110100110000" => B1 := "1011111"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3377
		when "110100110001" => B1 := "1110000"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3378
		when "110100110010" => B1 := "1111111"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3379
		when "110100110011" => B1 := "1111011"; B2 := "1110000"; B3 := "1111001"; B4 := "1111001"; 
		--3380
		when "110100110100" => B1 := "1111110"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3381
		when "110100110101" => B1 := "0110000"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3382
		when "110100110110" => B1 := "1101101"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3383
		when "110100110111" => B1 := "1111001"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3384
		when "110100111000" => B1 := "0110011"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3385
		when "110100111001" => B1 := "1011011"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3386
		when "110100111010" => B1 := "1011111"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3387
		when "110100111011" => B1 := "1110000"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3388
		when "110100111100" => B1 := "1111111"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3389
		when "110100111101" => B1 := "1111011"; B2 := "1111111"; B3 := "1111001"; B4 := "1111001"; 
		--3390
		when "110100111110" => B1 := "1111110"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3391
		when "110100111111" => B1 := "0110000"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3392
		when "110101000000" => B1 := "1101101"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3393
		when "110101000001" => B1 := "1111001"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3394
		when "110101000010" => B1 := "0110011"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3395
		when "110101000011" => B1 := "1011011"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3396
		when "110101000100" => B1 := "1011111"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3397
		when "110101000101" => B1 := "1110000"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3398
		when "110101000110" => B1 := "1111111"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3399
		when "110101000111" => B1 := "1111011"; B2 := "1111011"; B3 := "1111001"; B4 := "1111001"; 
		--3400
		when "110101001000" => B1 := "1111110"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3401
		when "110101001001" => B1 := "0110000"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3402
		when "110101001010" => B1 := "1101101"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3403
		when "110101001011" => B1 := "1111001"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3404
		when "110101001100" => B1 := "0110011"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3405
		when "110101001101" => B1 := "1011011"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3406
		when "110101001110" => B1 := "1011111"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3407
		when "110101001111" => B1 := "1110000"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3408
		when "110101010000" => B1 := "1111111"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3409
		when "110101010001" => B1 := "1111011"; B2 := "1111110"; B3 := "0110011"; B4 := "1111001"; 
		--3410
		when "110101010010" => B1 := "1111110"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3411
		when "110101010011" => B1 := "0110000"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3412
		when "110101010100" => B1 := "1101101"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3413
		when "110101010101" => B1 := "1111001"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3414
		when "110101010110" => B1 := "0110011"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3415
		when "110101010111" => B1 := "1011011"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3416
		when "110101011000" => B1 := "1011111"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3417
		when "110101011001" => B1 := "1110000"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3418
		when "110101011010" => B1 := "1111111"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3419
		when "110101011011" => B1 := "1111011"; B2 := "0110000"; B3 := "0110011"; B4 := "1111001"; 
		--3420
		when "110101011100" => B1 := "1111110"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3421
		when "110101011101" => B1 := "0110000"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3422
		when "110101011110" => B1 := "1101101"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3423
		when "110101011111" => B1 := "1111001"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3424
		when "110101100000" => B1 := "0110011"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3425
		when "110101100001" => B1 := "1011011"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3426
		when "110101100010" => B1 := "1011111"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3427
		when "110101100011" => B1 := "1110000"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3428
		when "110101100100" => B1 := "1111111"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3429
		when "110101100101" => B1 := "1111011"; B2 := "1101101"; B3 := "0110011"; B4 := "1111001"; 
		--3430
		when "110101100110" => B1 := "1111110"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3431
		when "110101100111" => B1 := "0110000"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3432
		when "110101101000" => B1 := "1101101"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3433
		when "110101101001" => B1 := "1111001"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3434
		when "110101101010" => B1 := "0110011"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3435
		when "110101101011" => B1 := "1011011"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3436
		when "110101101100" => B1 := "1011111"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3437
		when "110101101101" => B1 := "1110000"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3438
		when "110101101110" => B1 := "1111111"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3439
		when "110101101111" => B1 := "1111011"; B2 := "1111001"; B3 := "0110011"; B4 := "1111001"; 
		--3440
		when "110101110000" => B1 := "1111110"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3441
		when "110101110001" => B1 := "0110000"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3442
		when "110101110010" => B1 := "1101101"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3443
		when "110101110011" => B1 := "1111001"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3444
		when "110101110100" => B1 := "0110011"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3445
		when "110101110101" => B1 := "1011011"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3446
		when "110101110110" => B1 := "1011111"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3447
		when "110101110111" => B1 := "1110000"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3448
		when "110101111000" => B1 := "1111111"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3449
		when "110101111001" => B1 := "1111011"; B2 := "0110011"; B3 := "0110011"; B4 := "1111001"; 
		--3450
		when "110101111010" => B1 := "1111110"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3451
		when "110101111011" => B1 := "0110000"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3452
		when "110101111100" => B1 := "1101101"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3453
		when "110101111101" => B1 := "1111001"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3454
		when "110101111110" => B1 := "0110011"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3455
		when "110101111111" => B1 := "1011011"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3456
		when "110110000000" => B1 := "1011111"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3457
		when "110110000001" => B1 := "1110000"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3458
		when "110110000010" => B1 := "1111111"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3459
		when "110110000011" => B1 := "1111011"; B2 := "1011011"; B3 := "0110011"; B4 := "1111001"; 
		--3460
		when "110110000100" => B1 := "1111110"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3461
		when "110110000101" => B1 := "0110000"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3462
		when "110110000110" => B1 := "1101101"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3463
		when "110110000111" => B1 := "1111001"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3464
		when "110110001000" => B1 := "0110011"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3465
		when "110110001001" => B1 := "1011011"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3466
		when "110110001010" => B1 := "1011111"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3467
		when "110110001011" => B1 := "1110000"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3468
		when "110110001100" => B1 := "1111111"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3469
		when "110110001101" => B1 := "1111011"; B2 := "1011111"; B3 := "0110011"; B4 := "1111001"; 
		--3470
		when "110110001110" => B1 := "1111110"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3471
		when "110110001111" => B1 := "0110000"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3472
		when "110110010000" => B1 := "1101101"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3473
		when "110110010001" => B1 := "1111001"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3474
		when "110110010010" => B1 := "0110011"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3475
		when "110110010011" => B1 := "1011011"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3476
		when "110110010100" => B1 := "1011111"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3477
		when "110110010101" => B1 := "1110000"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3478
		when "110110010110" => B1 := "1111111"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3479
		when "110110010111" => B1 := "1111011"; B2 := "1110000"; B3 := "0110011"; B4 := "1111001"; 
		--3480
		when "110110011000" => B1 := "1111110"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3481
		when "110110011001" => B1 := "0110000"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3482
		when "110110011010" => B1 := "1101101"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3483
		when "110110011011" => B1 := "1111001"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3484
		when "110110011100" => B1 := "0110011"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3485
		when "110110011101" => B1 := "1011011"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3486
		when "110110011110" => B1 := "1011111"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3487
		when "110110011111" => B1 := "1110000"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3488
		when "110110100000" => B1 := "1111111"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3489
		when "110110100001" => B1 := "1111011"; B2 := "1111111"; B3 := "0110011"; B4 := "1111001"; 
		--3490
		when "110110100010" => B1 := "1111110"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3491
		when "110110100011" => B1 := "0110000"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3492
		when "110110100100" => B1 := "1101101"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3493
		when "110110100101" => B1 := "1111001"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3494
		when "110110100110" => B1 := "0110011"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3495
		when "110110100111" => B1 := "1011011"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3496
		when "110110101000" => B1 := "1011111"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3497
		when "110110101001" => B1 := "1110000"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3498
		when "110110101010" => B1 := "1111111"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3499
		when "110110101011" => B1 := "1111011"; B2 := "1111011"; B3 := "0110011"; B4 := "1111001"; 
		--3500
		when "110110101100" => B1 := "1111110"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3501
		when "110110101101" => B1 := "0110000"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3502
		when "110110101110" => B1 := "1101101"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3503
		when "110110101111" => B1 := "1111001"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3504
		when "110110110000" => B1 := "0110011"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3505
		when "110110110001" => B1 := "1011011"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3506
		when "110110110010" => B1 := "1011111"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3507
		when "110110110011" => B1 := "1110000"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3508
		when "110110110100" => B1 := "1111111"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3509
		when "110110110101" => B1 := "1111011"; B2 := "1111110"; B3 := "1011011"; B4 := "1111001"; 
		--3510
		when "110110110110" => B1 := "1111110"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3511
		when "110110110111" => B1 := "0110000"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3512
		when "110110111000" => B1 := "1101101"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3513
		when "110110111001" => B1 := "1111001"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3514
		when "110110111010" => B1 := "0110011"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3515
		when "110110111011" => B1 := "1011011"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3516
		when "110110111100" => B1 := "1011111"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3517
		when "110110111101" => B1 := "1110000"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3518
		when "110110111110" => B1 := "1111111"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3519
		when "110110111111" => B1 := "1111011"; B2 := "0110000"; B3 := "1011011"; B4 := "1111001"; 
		--3520
		when "110111000000" => B1 := "1111110"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3521
		when "110111000001" => B1 := "0110000"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3522
		when "110111000010" => B1 := "1101101"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3523
		when "110111000011" => B1 := "1111001"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3524
		when "110111000100" => B1 := "0110011"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3525
		when "110111000101" => B1 := "1011011"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3526
		when "110111000110" => B1 := "1011111"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3527
		when "110111000111" => B1 := "1110000"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3528
		when "110111001000" => B1 := "1111111"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3529
		when "110111001001" => B1 := "1111011"; B2 := "1101101"; B3 := "1011011"; B4 := "1111001"; 
		--3530
		when "110111001010" => B1 := "1111110"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3531
		when "110111001011" => B1 := "0110000"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3532
		when "110111001100" => B1 := "1101101"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3533
		when "110111001101" => B1 := "1111001"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3534
		when "110111001110" => B1 := "0110011"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3535
		when "110111001111" => B1 := "1011011"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3536
		when "110111010000" => B1 := "1011111"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3537
		when "110111010001" => B1 := "1110000"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3538
		when "110111010010" => B1 := "1111111"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3539
		when "110111010011" => B1 := "1111011"; B2 := "1111001"; B3 := "1011011"; B4 := "1111001"; 
		--3540
		when "110111010100" => B1 := "1111110"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3541
		when "110111010101" => B1 := "0110000"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3542
		when "110111010110" => B1 := "1101101"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3543
		when "110111010111" => B1 := "1111001"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3544
		when "110111011000" => B1 := "0110011"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3545
		when "110111011001" => B1 := "1011011"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3546
		when "110111011010" => B1 := "1011111"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3547
		when "110111011011" => B1 := "1110000"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3548
		when "110111011100" => B1 := "1111111"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3549
		when "110111011101" => B1 := "1111011"; B2 := "0110011"; B3 := "1011011"; B4 := "1111001"; 
		--3550
		when "110111011110" => B1 := "1111110"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3551
		when "110111011111" => B1 := "0110000"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3552
		when "110111100000" => B1 := "1101101"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3553
		when "110111100001" => B1 := "1111001"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3554
		when "110111100010" => B1 := "0110011"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3555
		when "110111100011" => B1 := "1011011"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3556
		when "110111100100" => B1 := "1011111"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3557
		when "110111100101" => B1 := "1110000"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3558
		when "110111100110" => B1 := "1111111"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3559
		when "110111100111" => B1 := "1111011"; B2 := "1011011"; B3 := "1011011"; B4 := "1111001"; 
		--3560
		when "110111101000" => B1 := "1111110"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3561
		when "110111101001" => B1 := "0110000"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3562
		when "110111101010" => B1 := "1101101"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3563
		when "110111101011" => B1 := "1111001"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3564
		when "110111101100" => B1 := "0110011"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3565
		when "110111101101" => B1 := "1011011"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3566
		when "110111101110" => B1 := "1011111"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3567
		when "110111101111" => B1 := "1110000"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3568
		when "110111110000" => B1 := "1111111"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3569
		when "110111110001" => B1 := "1111011"; B2 := "1011111"; B3 := "1011011"; B4 := "1111001"; 
		--3570
		when "110111110010" => B1 := "1111110"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3571
		when "110111110011" => B1 := "0110000"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3572
		when "110111110100" => B1 := "1101101"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3573
		when "110111110101" => B1 := "1111001"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3574
		when "110111110110" => B1 := "0110011"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3575
		when "110111110111" => B1 := "1011011"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3576
		when "110111111000" => B1 := "1011111"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3577
		when "110111111001" => B1 := "1110000"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3578
		when "110111111010" => B1 := "1111111"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3579
		when "110111111011" => B1 := "1111011"; B2 := "1110000"; B3 := "1011011"; B4 := "1111001"; 
		--3580
		when "110111111100" => B1 := "1111110"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3581
		when "110111111101" => B1 := "0110000"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3582
		when "110111111110" => B1 := "1101101"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3583
		when "110111111111" => B1 := "1111001"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3584
		when "111000000000" => B1 := "0110011"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3585
		when "111000000001" => B1 := "1011011"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3586
		when "111000000010" => B1 := "1011111"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3587
		when "111000000011" => B1 := "1110000"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3588
		when "111000000100" => B1 := "1111111"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3589
		when "111000000101" => B1 := "1111011"; B2 := "1111111"; B3 := "1011011"; B4 := "1111001"; 
		--3590
		when "111000000110" => B1 := "1111110"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3591
		when "111000000111" => B1 := "0110000"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3592
		when "111000001000" => B1 := "1101101"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3593
		when "111000001001" => B1 := "1111001"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3594
		when "111000001010" => B1 := "0110011"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3595
		when "111000001011" => B1 := "1011011"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3596
		when "111000001100" => B1 := "1011111"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3597
		when "111000001101" => B1 := "1110000"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3598
		when "111000001110" => B1 := "1111111"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3599
		when "111000001111" => B1 := "1111011"; B2 := "1111011"; B3 := "1011011"; B4 := "1111001"; 
		--3600
		when "111000010000" => B1 := "1111110"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3601
		when "111000010001" => B1 := "0110000"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3602
		when "111000010010" => B1 := "1101101"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3603
		when "111000010011" => B1 := "1111001"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3604
		when "111000010100" => B1 := "0110011"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3605
		when "111000010101" => B1 := "1011011"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3606
		when "111000010110" => B1 := "1011111"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3607
		when "111000010111" => B1 := "1110000"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3608
		when "111000011000" => B1 := "1111111"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3609
		when "111000011001" => B1 := "1111011"; B2 := "1111110"; B3 := "1011111"; B4 := "1111001"; 
		--3610
		when "111000011010" => B1 := "1111110"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3611
		when "111000011011" => B1 := "0110000"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3612
		when "111000011100" => B1 := "1101101"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3613
		when "111000011101" => B1 := "1111001"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3614
		when "111000011110" => B1 := "0110011"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3615
		when "111000011111" => B1 := "1011011"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3616
		when "111000100000" => B1 := "1011111"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3617
		when "111000100001" => B1 := "1110000"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3618
		when "111000100010" => B1 := "1111111"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3619
		when "111000100011" => B1 := "1111011"; B2 := "0110000"; B3 := "1011111"; B4 := "1111001"; 
		--3620
		when "111000100100" => B1 := "1111110"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3621
		when "111000100101" => B1 := "0110000"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3622
		when "111000100110" => B1 := "1101101"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3623
		when "111000100111" => B1 := "1111001"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3624
		when "111000101000" => B1 := "0110011"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3625
		when "111000101001" => B1 := "1011011"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3626
		when "111000101010" => B1 := "1011111"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3627
		when "111000101011" => B1 := "1110000"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3628
		when "111000101100" => B1 := "1111111"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3629
		when "111000101101" => B1 := "1111011"; B2 := "1101101"; B3 := "1011111"; B4 := "1111001"; 
		--3630
		when "111000101110" => B1 := "1111110"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3631
		when "111000101111" => B1 := "0110000"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3632
		when "111000110000" => B1 := "1101101"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3633
		when "111000110001" => B1 := "1111001"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3634
		when "111000110010" => B1 := "0110011"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3635
		when "111000110011" => B1 := "1011011"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3636
		when "111000110100" => B1 := "1011111"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3637
		when "111000110101" => B1 := "1110000"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3638
		when "111000110110" => B1 := "1111111"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3639
		when "111000110111" => B1 := "1111011"; B2 := "1111001"; B3 := "1011111"; B4 := "1111001"; 
		--3640
		when "111000111000" => B1 := "1111110"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3641
		when "111000111001" => B1 := "0110000"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3642
		when "111000111010" => B1 := "1101101"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3643
		when "111000111011" => B1 := "1111001"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3644
		when "111000111100" => B1 := "0110011"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3645
		when "111000111101" => B1 := "1011011"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3646
		when "111000111110" => B1 := "1011111"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3647
		when "111000111111" => B1 := "1110000"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3648
		when "111001000000" => B1 := "1111111"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3649
		when "111001000001" => B1 := "1111011"; B2 := "0110011"; B3 := "1011111"; B4 := "1111001"; 
		--3650
		when "111001000010" => B1 := "1111110"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3651
		when "111001000011" => B1 := "0110000"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3652
		when "111001000100" => B1 := "1101101"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3653
		when "111001000101" => B1 := "1111001"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3654
		when "111001000110" => B1 := "0110011"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3655
		when "111001000111" => B1 := "1011011"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3656
		when "111001001000" => B1 := "1011111"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3657
		when "111001001001" => B1 := "1110000"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3658
		when "111001001010" => B1 := "1111111"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3659
		when "111001001011" => B1 := "1111011"; B2 := "1011011"; B3 := "1011111"; B4 := "1111001"; 
		--3660
		when "111001001100" => B1 := "1111110"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3661
		when "111001001101" => B1 := "0110000"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3662
		when "111001001110" => B1 := "1101101"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3663
		when "111001001111" => B1 := "1111001"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3664
		when "111001010000" => B1 := "0110011"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3665
		when "111001010001" => B1 := "1011011"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3666
		when "111001010010" => B1 := "1011111"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3667
		when "111001010011" => B1 := "1110000"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3668
		when "111001010100" => B1 := "1111111"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3669
		when "111001010101" => B1 := "1111011"; B2 := "1011111"; B3 := "1011111"; B4 := "1111001"; 
		--3670
		when "111001010110" => B1 := "1111110"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3671
		when "111001010111" => B1 := "0110000"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3672
		when "111001011000" => B1 := "1101101"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3673
		when "111001011001" => B1 := "1111001"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3674
		when "111001011010" => B1 := "0110011"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3675
		when "111001011011" => B1 := "1011011"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3676
		when "111001011100" => B1 := "1011111"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3677
		when "111001011101" => B1 := "1110000"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3678
		when "111001011110" => B1 := "1111111"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3679
		when "111001011111" => B1 := "1111011"; B2 := "1110000"; B3 := "1011111"; B4 := "1111001"; 
		--3680
		when "111001100000" => B1 := "1111110"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3681
		when "111001100001" => B1 := "0110000"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3682
		when "111001100010" => B1 := "1101101"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3683
		when "111001100011" => B1 := "1111001"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3684
		when "111001100100" => B1 := "0110011"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3685
		when "111001100101" => B1 := "1011011"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3686
		when "111001100110" => B1 := "1011111"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3687
		when "111001100111" => B1 := "1110000"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3688
		when "111001101000" => B1 := "1111111"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3689
		when "111001101001" => B1 := "1111011"; B2 := "1111111"; B3 := "1011111"; B4 := "1111001"; 
		--3690
		when "111001101010" => B1 := "1111110"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3691
		when "111001101011" => B1 := "0110000"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3692
		when "111001101100" => B1 := "1101101"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3693
		when "111001101101" => B1 := "1111001"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3694
		when "111001101110" => B1 := "0110011"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3695
		when "111001101111" => B1 := "1011011"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3696
		when "111001110000" => B1 := "1011111"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3697
		when "111001110001" => B1 := "1110000"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3698
		when "111001110010" => B1 := "1111111"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3699
		when "111001110011" => B1 := "1111011"; B2 := "1111011"; B3 := "1011111"; B4 := "1111001"; 
		--3700
		when "111001110100" => B1 := "1111110"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3701
		when "111001110101" => B1 := "0110000"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3702
		when "111001110110" => B1 := "1101101"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3703
		when "111001110111" => B1 := "1111001"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3704
		when "111001111000" => B1 := "0110011"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3705
		when "111001111001" => B1 := "1011011"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3706
		when "111001111010" => B1 := "1011111"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3707
		when "111001111011" => B1 := "1110000"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3708
		when "111001111100" => B1 := "1111111"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3709
		when "111001111101" => B1 := "1111011"; B2 := "1111110"; B3 := "1110000"; B4 := "1111001"; 
		--3710
		when "111001111110" => B1 := "1111110"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3711
		when "111001111111" => B1 := "0110000"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3712
		when "111010000000" => B1 := "1101101"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3713
		when "111010000001" => B1 := "1111001"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3714
		when "111010000010" => B1 := "0110011"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3715
		when "111010000011" => B1 := "1011011"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3716
		when "111010000100" => B1 := "1011111"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3717
		when "111010000101" => B1 := "1110000"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3718
		when "111010000110" => B1 := "1111111"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3719
		when "111010000111" => B1 := "1111011"; B2 := "0110000"; B3 := "1110000"; B4 := "1111001"; 
		--3720
		when "111010001000" => B1 := "1111110"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3721
		when "111010001001" => B1 := "0110000"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3722
		when "111010001010" => B1 := "1101101"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3723
		when "111010001011" => B1 := "1111001"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3724
		when "111010001100" => B1 := "0110011"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3725
		when "111010001101" => B1 := "1011011"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3726
		when "111010001110" => B1 := "1011111"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3727
		when "111010001111" => B1 := "1110000"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3728
		when "111010010000" => B1 := "1111111"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3729
		when "111010010001" => B1 := "1111011"; B2 := "1101101"; B3 := "1110000"; B4 := "1111001"; 
		--3730
		when "111010010010" => B1 := "1111110"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3731
		when "111010010011" => B1 := "0110000"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3732
		when "111010010100" => B1 := "1101101"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3733
		when "111010010101" => B1 := "1111001"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3734
		when "111010010110" => B1 := "0110011"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3735
		when "111010010111" => B1 := "1011011"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3736
		when "111010011000" => B1 := "1011111"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3737
		when "111010011001" => B1 := "1110000"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3738
		when "111010011010" => B1 := "1111111"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3739
		when "111010011011" => B1 := "1111011"; B2 := "1111001"; B3 := "1110000"; B4 := "1111001"; 
		--3740
		when "111010011100" => B1 := "1111110"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3741
		when "111010011101" => B1 := "0110000"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3742
		when "111010011110" => B1 := "1101101"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3743
		when "111010011111" => B1 := "1111001"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3744
		when "111010100000" => B1 := "0110011"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3745
		when "111010100001" => B1 := "1011011"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3746
		when "111010100010" => B1 := "1011111"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3747
		when "111010100011" => B1 := "1110000"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3748
		when "111010100100" => B1 := "1111111"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3749
		when "111010100101" => B1 := "1111011"; B2 := "0110011"; B3 := "1110000"; B4 := "1111001"; 
		--3750
		when "111010100110" => B1 := "1111110"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3751
		when "111010100111" => B1 := "0110000"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3752
		when "111010101000" => B1 := "1101101"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3753
		when "111010101001" => B1 := "1111001"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3754
		when "111010101010" => B1 := "0110011"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3755
		when "111010101011" => B1 := "1011011"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3756
		when "111010101100" => B1 := "1011111"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3757
		when "111010101101" => B1 := "1110000"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3758
		when "111010101110" => B1 := "1111111"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3759
		when "111010101111" => B1 := "1111011"; B2 := "1011011"; B3 := "1110000"; B4 := "1111001"; 
		--3760
		when "111010110000" => B1 := "1111110"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3761
		when "111010110001" => B1 := "0110000"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3762
		when "111010110010" => B1 := "1101101"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3763
		when "111010110011" => B1 := "1111001"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3764
		when "111010110100" => B1 := "0110011"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3765
		when "111010110101" => B1 := "1011011"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3766
		when "111010110110" => B1 := "1011111"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3767
		when "111010110111" => B1 := "1110000"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3768
		when "111010111000" => B1 := "1111111"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3769
		when "111010111001" => B1 := "1111011"; B2 := "1011111"; B3 := "1110000"; B4 := "1111001"; 
		--3770
		when "111010111010" => B1 := "1111110"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3771
		when "111010111011" => B1 := "0110000"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3772
		when "111010111100" => B1 := "1101101"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3773
		when "111010111101" => B1 := "1111001"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3774
		when "111010111110" => B1 := "0110011"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3775
		when "111010111111" => B1 := "1011011"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3776
		when "111011000000" => B1 := "1011111"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3777
		when "111011000001" => B1 := "1110000"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3778
		when "111011000010" => B1 := "1111111"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3779
		when "111011000011" => B1 := "1111011"; B2 := "1110000"; B3 := "1110000"; B4 := "1111001"; 
		--3780
		when "111011000100" => B1 := "1111110"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3781
		when "111011000101" => B1 := "0110000"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3782
		when "111011000110" => B1 := "1101101"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3783
		when "111011000111" => B1 := "1111001"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3784
		when "111011001000" => B1 := "0110011"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3785
		when "111011001001" => B1 := "1011011"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3786
		when "111011001010" => B1 := "1011111"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3787
		when "111011001011" => B1 := "1110000"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3788
		when "111011001100" => B1 := "1111111"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3789
		when "111011001101" => B1 := "1111011"; B2 := "1111111"; B3 := "1110000"; B4 := "1111001"; 
		--3790
		when "111011001110" => B1 := "1111110"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3791
		when "111011001111" => B1 := "0110000"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3792
		when "111011010000" => B1 := "1101101"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3793
		when "111011010001" => B1 := "1111001"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3794
		when "111011010010" => B1 := "0110011"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3795
		when "111011010011" => B1 := "1011011"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3796
		when "111011010100" => B1 := "1011111"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3797
		when "111011010101" => B1 := "1110000"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3798
		when "111011010110" => B1 := "1111111"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3799
		when "111011010111" => B1 := "1111011"; B2 := "1111011"; B3 := "1110000"; B4 := "1111001"; 
		--3800
		when "111011011000" => B1 := "1111110"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3801
		when "111011011001" => B1 := "0110000"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3802
		when "111011011010" => B1 := "1101101"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3803
		when "111011011011" => B1 := "1111001"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3804
		when "111011011100" => B1 := "0110011"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3805
		when "111011011101" => B1 := "1011011"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3806
		when "111011011110" => B1 := "1011111"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3807
		when "111011011111" => B1 := "1110000"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3808
		when "111011100000" => B1 := "1111111"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3809
		when "111011100001" => B1 := "1111011"; B2 := "1111110"; B3 := "1111111"; B4 := "1111001"; 
		--3810
		when "111011100010" => B1 := "1111110"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3811
		when "111011100011" => B1 := "0110000"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3812
		when "111011100100" => B1 := "1101101"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3813
		when "111011100101" => B1 := "1111001"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3814
		when "111011100110" => B1 := "0110011"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3815
		when "111011100111" => B1 := "1011011"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3816
		when "111011101000" => B1 := "1011111"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3817
		when "111011101001" => B1 := "1110000"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3818
		when "111011101010" => B1 := "1111111"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3819
		when "111011101011" => B1 := "1111011"; B2 := "0110000"; B3 := "1111111"; B4 := "1111001"; 
		--3820
		when "111011101100" => B1 := "1111110"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3821
		when "111011101101" => B1 := "0110000"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3822
		when "111011101110" => B1 := "1101101"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3823
		when "111011101111" => B1 := "1111001"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3824
		when "111011110000" => B1 := "0110011"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3825
		when "111011110001" => B1 := "1011011"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3826
		when "111011110010" => B1 := "1011111"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3827
		when "111011110011" => B1 := "1110000"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3828
		when "111011110100" => B1 := "1111111"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3829
		when "111011110101" => B1 := "1111011"; B2 := "1101101"; B3 := "1111111"; B4 := "1111001"; 
		--3830
		when "111011110110" => B1 := "1111110"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3831
		when "111011110111" => B1 := "0110000"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3832
		when "111011111000" => B1 := "1101101"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3833
		when "111011111001" => B1 := "1111001"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3834
		when "111011111010" => B1 := "0110011"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3835
		when "111011111011" => B1 := "1011011"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3836
		when "111011111100" => B1 := "1011111"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3837
		when "111011111101" => B1 := "1110000"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3838
		when "111011111110" => B1 := "1111111"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3839
		when "111011111111" => B1 := "1111011"; B2 := "1111001"; B3 := "1111111"; B4 := "1111001"; 
		--3840
		when "111100000000" => B1 := "1111110"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3841
		when "111100000001" => B1 := "0110000"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3842
		when "111100000010" => B1 := "1101101"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3843
		when "111100000011" => B1 := "1111001"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3844
		when "111100000100" => B1 := "0110011"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3845
		when "111100000101" => B1 := "1011011"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3846
		when "111100000110" => B1 := "1011111"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3847
		when "111100000111" => B1 := "1110000"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3848
		when "111100001000" => B1 := "1111111"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3849
		when "111100001001" => B1 := "1111011"; B2 := "0110011"; B3 := "1111111"; B4 := "1111001"; 
		--3850
		when "111100001010" => B1 := "1111110"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3851
		when "111100001011" => B1 := "0110000"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3852
		when "111100001100" => B1 := "1101101"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3853
		when "111100001101" => B1 := "1111001"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3854
		when "111100001110" => B1 := "0110011"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3855
		when "111100001111" => B1 := "1011011"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3856
		when "111100010000" => B1 := "1011111"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3857
		when "111100010001" => B1 := "1110000"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3858
		when "111100010010" => B1 := "1111111"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3859
		when "111100010011" => B1 := "1111011"; B2 := "1011011"; B3 := "1111111"; B4 := "1111001"; 
		--3860
		when "111100010100" => B1 := "1111110"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3861
		when "111100010101" => B1 := "0110000"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3862
		when "111100010110" => B1 := "1101101"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3863
		when "111100010111" => B1 := "1111001"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3864
		when "111100011000" => B1 := "0110011"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3865
		when "111100011001" => B1 := "1011011"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3866
		when "111100011010" => B1 := "1011111"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3867
		when "111100011011" => B1 := "1110000"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3868
		when "111100011100" => B1 := "1111111"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3869
		when "111100011101" => B1 := "1111011"; B2 := "1011111"; B3 := "1111111"; B4 := "1111001"; 
		--3870
		when "111100011110" => B1 := "1111110"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3871
		when "111100011111" => B1 := "0110000"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3872
		when "111100100000" => B1 := "1101101"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3873
		when "111100100001" => B1 := "1111001"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3874
		when "111100100010" => B1 := "0110011"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3875
		when "111100100011" => B1 := "1011011"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3876
		when "111100100100" => B1 := "1011111"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3877
		when "111100100101" => B1 := "1110000"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3878
		when "111100100110" => B1 := "1111111"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3879
		when "111100100111" => B1 := "1111011"; B2 := "1110000"; B3 := "1111111"; B4 := "1111001"; 
		--3880
		when "111100101000" => B1 := "1111110"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3881
		when "111100101001" => B1 := "0110000"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3882
		when "111100101010" => B1 := "1101101"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3883
		when "111100101011" => B1 := "1111001"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3884
		when "111100101100" => B1 := "0110011"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3885
		when "111100101101" => B1 := "1011011"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3886
		when "111100101110" => B1 := "1011111"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3887
		when "111100101111" => B1 := "1110000"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3888
		when "111100110000" => B1 := "1111111"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3889
		when "111100110001" => B1 := "1111011"; B2 := "1111111"; B3 := "1111111"; B4 := "1111001"; 
		--3890
		when "111100110010" => B1 := "1111110"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3891
		when "111100110011" => B1 := "0110000"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3892
		when "111100110100" => B1 := "1101101"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3893
		when "111100110101" => B1 := "1111001"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3894
		when "111100110110" => B1 := "0110011"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3895
		when "111100110111" => B1 := "1011011"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3896
		when "111100111000" => B1 := "1011111"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3897
		when "111100111001" => B1 := "1110000"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3898
		when "111100111010" => B1 := "1111111"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3899
		when "111100111011" => B1 := "1111011"; B2 := "1111011"; B3 := "1111111"; B4 := "1111001"; 
		--3900
		when "111100111100" => B1 := "1111110"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3901
		when "111100111101" => B1 := "0110000"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3902
		when "111100111110" => B1 := "1101101"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3903
		when "111100111111" => B1 := "1111001"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3904
		when "111101000000" => B1 := "0110011"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3905
		when "111101000001" => B1 := "1011011"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3906
		when "111101000010" => B1 := "1011111"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3907
		when "111101000011" => B1 := "1110000"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3908
		when "111101000100" => B1 := "1111111"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3909
		when "111101000101" => B1 := "1111011"; B2 := "1111110"; B3 := "1111011"; B4 := "1111001"; 
		--3910
		when "111101000110" => B1 := "1111110"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3911
		when "111101000111" => B1 := "0110000"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3912
		when "111101001000" => B1 := "1101101"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3913
		when "111101001001" => B1 := "1111001"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3914
		when "111101001010" => B1 := "0110011"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3915
		when "111101001011" => B1 := "1011011"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3916
		when "111101001100" => B1 := "1011111"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3917
		when "111101001101" => B1 := "1110000"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3918
		when "111101001110" => B1 := "1111111"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3919
		when "111101001111" => B1 := "1111011"; B2 := "0110000"; B3 := "1111011"; B4 := "1111001"; 
		--3920
		when "111101010000" => B1 := "1111110"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3921
		when "111101010001" => B1 := "0110000"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3922
		when "111101010010" => B1 := "1101101"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3923
		when "111101010011" => B1 := "1111001"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3924
		when "111101010100" => B1 := "0110011"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3925
		when "111101010101" => B1 := "1011011"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3926
		when "111101010110" => B1 := "1011111"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3927
		when "111101010111" => B1 := "1110000"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3928
		when "111101011000" => B1 := "1111111"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3929
		when "111101011001" => B1 := "1111011"; B2 := "1101101"; B3 := "1111011"; B4 := "1111001"; 
		--3930
		when "111101011010" => B1 := "1111110"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3931
		when "111101011011" => B1 := "0110000"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3932
		when "111101011100" => B1 := "1101101"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3933
		when "111101011101" => B1 := "1111001"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3934
		when "111101011110" => B1 := "0110011"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3935
		when "111101011111" => B1 := "1011011"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3936
		when "111101100000" => B1 := "1011111"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3937
		when "111101100001" => B1 := "1110000"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3938
		when "111101100010" => B1 := "1111111"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3939
		when "111101100011" => B1 := "1111011"; B2 := "1111001"; B3 := "1111011"; B4 := "1111001"; 
		--3940
		when "111101100100" => B1 := "1111110"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3941
		when "111101100101" => B1 := "0110000"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3942
		when "111101100110" => B1 := "1101101"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3943
		when "111101100111" => B1 := "1111001"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3944
		when "111101101000" => B1 := "0110011"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3945
		when "111101101001" => B1 := "1011011"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3946
		when "111101101010" => B1 := "1011111"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3947
		when "111101101011" => B1 := "1110000"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3948
		when "111101101100" => B1 := "1111111"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3949
		when "111101101101" => B1 := "1111011"; B2 := "0110011"; B3 := "1111011"; B4 := "1111001"; 
		--3950
		when "111101101110" => B1 := "1111110"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3951
		when "111101101111" => B1 := "0110000"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3952
		when "111101110000" => B1 := "1101101"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3953
		when "111101110001" => B1 := "1111001"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3954
		when "111101110010" => B1 := "0110011"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3955
		when "111101110011" => B1 := "1011011"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3956
		when "111101110100" => B1 := "1011111"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3957
		when "111101110101" => B1 := "1110000"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3958
		when "111101110110" => B1 := "1111111"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3959
		when "111101110111" => B1 := "1111011"; B2 := "1011011"; B3 := "1111011"; B4 := "1111001"; 
		--3960
		when "111101111000" => B1 := "1111110"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3961
		when "111101111001" => B1 := "0110000"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3962
		when "111101111010" => B1 := "1101101"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3963
		when "111101111011" => B1 := "1111001"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3964
		when "111101111100" => B1 := "0110011"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3965
		when "111101111101" => B1 := "1011011"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3966
		when "111101111110" => B1 := "1011111"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3967
		when "111101111111" => B1 := "1110000"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3968
		when "111110000000" => B1 := "1111111"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3969
		when "111110000001" => B1 := "1111011"; B2 := "1011111"; B3 := "1111011"; B4 := "1111001"; 
		--3970
		when "111110000010" => B1 := "1111110"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3971
		when "111110000011" => B1 := "0110000"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3972
		when "111110000100" => B1 := "1101101"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3973
		when "111110000101" => B1 := "1111001"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3974
		when "111110000110" => B1 := "0110011"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3975
		when "111110000111" => B1 := "1011011"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3976
		when "111110001000" => B1 := "1011111"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3977
		when "111110001001" => B1 := "1110000"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3978
		when "111110001010" => B1 := "1111111"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3979
		when "111110001011" => B1 := "1111011"; B2 := "1110000"; B3 := "1111011"; B4 := "1111001"; 
		--3980
		when "111110001100" => B1 := "1111110"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3981
		when "111110001101" => B1 := "0110000"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3982
		when "111110001110" => B1 := "1101101"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3983
		when "111110001111" => B1 := "1111001"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3984
		when "111110010000" => B1 := "0110011"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3985
		when "111110010001" => B1 := "1011011"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3986
		when "111110010010" => B1 := "1011111"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3987
		when "111110010011" => B1 := "1110000"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3988
		when "111110010100" => B1 := "1111111"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3989
		when "111110010101" => B1 := "1111011"; B2 := "1111111"; B3 := "1111011"; B4 := "1111001"; 
		--3990
		when "111110010110" => B1 := "1111110"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--3991
		when "111110010111" => B1 := "0110000"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--3992
		when "111110011000" => B1 := "1101101"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--3993
		when "111110011001" => B1 := "1111001"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--3994
		when "111110011010" => B1 := "0110011"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--3995
		when "111110011011" => B1 := "1011011"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--3996
		when "111110011100" => B1 := "1011111"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--3997
		when "111110011101" => B1 := "1110000"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--3998
		when "111110011110" => B1 := "1111111"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--3999
		when "111110011111" => B1 := "1111011"; B2 := "1111011"; B3 := "1111011"; B4 := "1111001"; 
		--4000
		when "111110100000" => B1 := "1111110"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4001
		when "111110100001" => B1 := "0110000"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4002
		when "111110100010" => B1 := "1101101"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4003
		when "111110100011" => B1 := "1111001"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4004
		when "111110100100" => B1 := "0110011"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4005
		when "111110100101" => B1 := "1011011"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4006
		when "111110100110" => B1 := "1011111"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4007
		when "111110100111" => B1 := "1110000"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4008
		when "111110101000" => B1 := "1111111"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4009
		when "111110101001" => B1 := "1111011"; B2 := "1111110"; B3 := "1111110"; B4 := "0110011"; 
		--4010
		when "111110101010" => B1 := "1111110"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4011
		when "111110101011" => B1 := "0110000"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4012
		when "111110101100" => B1 := "1101101"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4013
		when "111110101101" => B1 := "1111001"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4014
		when "111110101110" => B1 := "0110011"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4015
		when "111110101111" => B1 := "1011011"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4016
		when "111110110000" => B1 := "1011111"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4017
		when "111110110001" => B1 := "1110000"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4018
		when "111110110010" => B1 := "1111111"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4019
		when "111110110011" => B1 := "1111011"; B2 := "0110000"; B3 := "1111110"; B4 := "0110011"; 
		--4020
		when "111110110100" => B1 := "1111110"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4021
		when "111110110101" => B1 := "0110000"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4022
		when "111110110110" => B1 := "1101101"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4023
		when "111110110111" => B1 := "1111001"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4024
		when "111110111000" => B1 := "0110011"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4025
		when "111110111001" => B1 := "1011011"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4026
		when "111110111010" => B1 := "1011111"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4027
		when "111110111011" => B1 := "1110000"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4028
		when "111110111100" => B1 := "1111111"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4029
		when "111110111101" => B1 := "1111011"; B2 := "1101101"; B3 := "1111110"; B4 := "0110011"; 
		--4030
		when "111110111110" => B1 := "1111110"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4031
		when "111110111111" => B1 := "0110000"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4032
		when "111111000000" => B1 := "1101101"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4033
		when "111111000001" => B1 := "1111001"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4034
		when "111111000010" => B1 := "0110011"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4035
		when "111111000011" => B1 := "1011011"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4036
		when "111111000100" => B1 := "1011111"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4037
		when "111111000101" => B1 := "1110000"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4038
		when "111111000110" => B1 := "1111111"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4039
		when "111111000111" => B1 := "1111011"; B2 := "1111001"; B3 := "1111110"; B4 := "0110011"; 
		--4040
		when "111111001000" => B1 := "1111110"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4041
		when "111111001001" => B1 := "0110000"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4042
		when "111111001010" => B1 := "1101101"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4043
		when "111111001011" => B1 := "1111001"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4044
		when "111111001100" => B1 := "0110011"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4045
		when "111111001101" => B1 := "1011011"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4046
		when "111111001110" => B1 := "1011111"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4047
		when "111111001111" => B1 := "1110000"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4048
		when "111111010000" => B1 := "1111111"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4049
		when "111111010001" => B1 := "1111011"; B2 := "0110011"; B3 := "1111110"; B4 := "0110011"; 
		--4050
		when "111111010010" => B1 := "1111110"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4051
		when "111111010011" => B1 := "0110000"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4052
		when "111111010100" => B1 := "1101101"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4053
		when "111111010101" => B1 := "1111001"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4054
		when "111111010110" => B1 := "0110011"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4055
		when "111111010111" => B1 := "1011011"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4056
		when "111111011000" => B1 := "1011111"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4057
		when "111111011001" => B1 := "1110000"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4058
		when "111111011010" => B1 := "1111111"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4059
		when "111111011011" => B1 := "1111011"; B2 := "1011011"; B3 := "1111110"; B4 := "0110011"; 
		--4060
		when "111111011100" => B1 := "1111110"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4061
		when "111111011101" => B1 := "0110000"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4062
		when "111111011110" => B1 := "1101101"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4063
		when "111111011111" => B1 := "1111001"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4064
		when "111111100000" => B1 := "0110011"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4065
		when "111111100001" => B1 := "1011011"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4066
		when "111111100010" => B1 := "1011111"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4067
		when "111111100011" => B1 := "1110000"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4068
		when "111111100100" => B1 := "1111111"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4069
		when "111111100101" => B1 := "1111011"; B2 := "1011111"; B3 := "1111110"; B4 := "0110011"; 
		--4070
		when "111111100110" => B1 := "1111110"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4071
		when "111111100111" => B1 := "0110000"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4072
		when "111111101000" => B1 := "1101101"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4073
		when "111111101001" => B1 := "1111001"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4074
		when "111111101010" => B1 := "0110011"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4075
		when "111111101011" => B1 := "1011011"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4076
		when "111111101100" => B1 := "1011111"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4077
		when "111111101101" => B1 := "1110000"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4078
		when "111111101110" => B1 := "1111111"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4079
		when "111111101111" => B1 := "1111011"; B2 := "1110000"; B3 := "1111110"; B4 := "0110011"; 
		--4080
		when "111111110000" => B1 := "1111110"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4081
		when "111111110001" => B1 := "0110000"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4082
		when "111111110010" => B1 := "1101101"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4083
		when "111111110011" => B1 := "1111001"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4084
		when "111111110100" => B1 := "0110011"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4085
		when "111111110101" => B1 := "1011011"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4086
		when "111111110110" => B1 := "1011111"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4087
		when "111111110111" => B1 := "1110000"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4088
		when "111111111000" => B1 := "1111111"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4089
		when "111111111001" => B1 := "1111011"; B2 := "1111111"; B3 := "1111110"; B4 := "0110011"; 
		--4090
		when "111111111010" => B1 := "1111110"; B2 := "1111011"; B3 := "1111110"; B4 := "0110011"; 
		--4091
		when "111111111011" => B1 := "0110000"; B2 := "1111011"; B3 := "1111110"; B4 := "0110011"; 
		--4092
		when "111111111100" => B1 := "1101101"; B2 := "1111011"; B3 := "1111110"; B4 := "0110011"; 
		--4093
		when "111111111101" => B1 := "1111001"; B2 := "1111011"; B3 := "1111110"; B4 := "0110011"; 
		--4094
		when "111111111110" => B1 := "0110011"; B2 := "1111011"; B3 := "1111110"; B4 := "0110011"; 
		--4095
		when "111111111111" => B1 := "1011011"; B2 := "1111011"; B3 := "1111110"; B4 := "0110011"; 

		when others => B1 := "XXXXXXX"; B2 := "XXXXXXX"; B3 := "XXXXXXX"; B4 := "XXXXXXX";
			
		end case;
		
		NRU<=B1;
		NRZ<=B2;
		NRS<=B3;
		NRM<=B4;
	
	end process;
	
end architecture;